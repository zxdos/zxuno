-------------------------------------------------------------------------------
--
-- Synthesizable model of TI's TMS9918A, TMS9928A, TMS9929A.
--
-- $Id: vdp18_col_mux-c.vhd,v 1.3 2006/06/18 10:47:01 arnim Exp $
--
-------------------------------------------------------------------------------

configuration vdp18_col_mux_rtl_c0 of vdp18_col_mux is

  for rtl
  end for;

end vdp18_col_mux_rtl_c0;
