
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity os8 is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(7 downto 0)
);
end os8;

architecture syn of os8 is
        type rom_type is array(0 to 8191) of std_logic_vector(7 downto 0);
        signal ROM:rom_type:=
(
	X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"18",
X"18",
X"00",
X"18",
X"00",
X"00",
X"66",
X"66",
X"66",
X"00",
X"00",
X"00",
X"00",
X"00",
X"66",
X"ff",
X"66",
X"66",
X"ff",
X"66",
X"00",
X"18",
X"3e",
X"60",
X"3c",
X"06",
X"7c",
X"18",
X"00",
X"00",
X"66",
X"6c",
X"18",
X"30",
X"66",
X"46",
X"00",
X"1c",
X"36",
X"1c",
X"38",
X"6f",
X"66",
X"3b",
X"00",
X"00",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"00",
X"00",
X"0e",
X"1c",
X"18",
X"18",
X"1c",
X"0e",
X"00",
X"00",
X"70",
X"38",
X"18",
X"18",
X"38",
X"70",
X"00",
X"00",
X"66",
X"3c",
X"ff",
X"3c",
X"66",
X"00",
X"00",
X"00",
X"18",
X"18",
X"7e",
X"18",
X"18",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"30",
X"00",
X"00",
X"00",
X"7e",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"00",
X"00",
X"06",
X"0c",
X"18",
X"30",
X"60",
X"40",
X"00",
X"00",
X"3c",
X"66",
X"6e",
X"76",
X"66",
X"3c",
X"00",
X"00",
X"18",
X"38",
X"18",
X"18",
X"18",
X"7e",
X"00",
X"00",
X"3c",
X"66",
X"0c",
X"18",
X"30",
X"7e",
X"00",
X"00",
X"7e",
X"0c",
X"18",
X"0c",
X"66",
X"3c",
X"00",
X"00",
X"0c",
X"1c",
X"3c",
X"6c",
X"7e",
X"0c",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"06",
X"66",
X"3c",
X"00",
X"00",
X"3c",
X"60",
X"7c",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"7e",
X"06",
X"0c",
X"18",
X"30",
X"30",
X"00",
X"00",
X"3c",
X"66",
X"3c",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"3c",
X"66",
X"3e",
X"06",
X"0c",
X"38",
X"00",
X"00",
X"00",
X"18",
X"18",
X"00",
X"18",
X"18",
X"00",
X"00",
X"00",
X"18",
X"18",
X"00",
X"18",
X"18",
X"30",
X"06",
X"0c",
X"18",
X"30",
X"18",
X"0c",
X"06",
X"00",
X"00",
X"00",
X"7e",
X"00",
X"00",
X"7e",
X"00",
X"00",
X"60",
X"30",
X"18",
X"0c",
X"18",
X"30",
X"60",
X"00",
X"00",
X"3c",
X"66",
X"0c",
X"18",
X"00",
X"18",
X"00",
X"00",
X"3c",
X"66",
X"6e",
X"6e",
X"60",
X"3e",
X"00",
X"00",
X"18",
X"3c",
X"66",
X"66",
X"7e",
X"66",
X"00",
X"00",
X"7c",
X"66",
X"7c",
X"66",
X"66",
X"7c",
X"00",
X"00",
X"3c",
X"66",
X"60",
X"60",
X"66",
X"3c",
X"00",
X"00",
X"78",
X"6c",
X"66",
X"66",
X"6c",
X"78",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"60",
X"60",
X"7e",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"60",
X"60",
X"60",
X"00",
X"00",
X"3e",
X"60",
X"60",
X"6e",
X"66",
X"3e",
X"00",
X"00",
X"66",
X"66",
X"7e",
X"66",
X"66",
X"66",
X"00",
X"00",
X"7e",
X"18",
X"18",
X"18",
X"18",
X"7e",
X"00",
X"00",
X"06",
X"06",
X"06",
X"06",
X"66",
X"3c",
X"00",
X"00",
X"66",
X"6c",
X"78",
X"78",
X"6c",
X"66",
X"00",
X"00",
X"60",
X"60",
X"60",
X"60",
X"60",
X"7e",
X"00",
X"00",
X"63",
X"77",
X"7f",
X"6b",
X"63",
X"63",
X"00",
X"00",
X"66",
X"76",
X"7e",
X"7e",
X"6e",
X"66",
X"00",
X"00",
X"3c",
X"66",
X"66",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"7c",
X"60",
X"60",
X"00",
X"00",
X"3c",
X"66",
X"66",
X"66",
X"6c",
X"36",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"7c",
X"6c",
X"66",
X"00",
X"00",
X"3c",
X"60",
X"3c",
X"06",
X"06",
X"3c",
X"00",
X"00",
X"7e",
X"18",
X"18",
X"18",
X"18",
X"18",
X"00",
X"00",
X"66",
X"66",
X"66",
X"66",
X"66",
X"7e",
X"00",
X"00",
X"66",
X"66",
X"66",
X"66",
X"3c",
X"18",
X"00",
X"00",
X"63",
X"63",
X"6b",
X"7f",
X"77",
X"63",
X"00",
X"00",
X"66",
X"66",
X"3c",
X"3c",
X"66",
X"66",
X"00",
X"00",
X"66",
X"66",
X"3c",
X"18",
X"18",
X"18",
X"00",
X"00",
X"7e",
X"0c",
X"18",
X"30",
X"60",
X"7e",
X"00",
X"00",
X"1e",
X"18",
X"18",
X"18",
X"18",
X"1e",
X"00",
X"00",
X"40",
X"60",
X"30",
X"18",
X"0c",
X"06",
X"00",
X"00",
X"78",
X"18",
X"18",
X"18",
X"18",
X"78",
X"00",
X"00",
X"08",
X"1c",
X"36",
X"63",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"00",
X"00",
X"36",
X"7f",
X"7f",
X"3e",
X"1c",
X"08",
X"00",
X"18",
X"18",
X"18",
X"1f",
X"1f",
X"18",
X"18",
X"18",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"18",
X"18",
X"18",
X"f8",
X"f8",
X"00",
X"00",
X"00",
X"18",
X"18",
X"18",
X"f8",
X"f8",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"f8",
X"f8",
X"18",
X"18",
X"18",
X"03",
X"07",
X"0e",
X"1c",
X"38",
X"70",
X"e0",
X"c0",
X"c0",
X"e0",
X"70",
X"38",
X"1c",
X"0e",
X"07",
X"03",
X"01",
X"03",
X"07",
X"0f",
X"1f",
X"3f",
X"7f",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"0f",
X"0f",
X"0f",
X"0f",
X"80",
X"c0",
X"e0",
X"f0",
X"f8",
X"fc",
X"fe",
X"ff",
X"0f",
X"0f",
X"0f",
X"0f",
X"00",
X"00",
X"00",
X"00",
X"f0",
X"f0",
X"f0",
X"f0",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"f0",
X"f0",
X"f0",
X"f0",
X"00",
X"1c",
X"1c",
X"77",
X"77",
X"08",
X"1c",
X"00",
X"00",
X"00",
X"00",
X"1f",
X"1f",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"18",
X"18",
X"18",
X"ff",
X"ff",
X"18",
X"18",
X"18",
X"00",
X"00",
X"3c",
X"7e",
X"7e",
X"7e",
X"3c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"c0",
X"c0",
X"c0",
X"c0",
X"c0",
X"c0",
X"c0",
X"c0",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"18",
X"18",
X"18",
X"1f",
X"1f",
X"00",
X"00",
X"00",
X"78",
X"60",
X"78",
X"60",
X"7e",
X"18",
X"1e",
X"00",
X"00",
X"18",
X"3c",
X"7e",
X"18",
X"18",
X"18",
X"00",
X"00",
X"18",
X"18",
X"18",
X"7e",
X"3c",
X"18",
X"00",
X"00",
X"18",
X"30",
X"7e",
X"30",
X"18",
X"00",
X"00",
X"00",
X"18",
X"0c",
X"7e",
X"0c",
X"18",
X"00",
X"00",
X"00",
X"18",
X"3c",
X"7e",
X"7e",
X"3c",
X"18",
X"00",
X"00",
X"00",
X"3c",
X"06",
X"3e",
X"66",
X"3e",
X"00",
X"00",
X"60",
X"60",
X"7c",
X"66",
X"66",
X"7c",
X"00",
X"00",
X"00",
X"3c",
X"60",
X"60",
X"60",
X"3c",
X"00",
X"00",
X"06",
X"06",
X"3e",
X"66",
X"66",
X"3e",
X"00",
X"00",
X"00",
X"3c",
X"66",
X"7e",
X"60",
X"3c",
X"00",
X"00",
X"0e",
X"18",
X"3e",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"3e",
X"66",
X"66",
X"3e",
X"06",
X"7c",
X"00",
X"60",
X"60",
X"7c",
X"66",
X"66",
X"66",
X"00",
X"00",
X"18",
X"00",
X"38",
X"18",
X"18",
X"3c",
X"00",
X"00",
X"06",
X"00",
X"06",
X"06",
X"06",
X"06",
X"3c",
X"00",
X"60",
X"60",
X"6c",
X"78",
X"6c",
X"66",
X"00",
X"00",
X"38",
X"18",
X"18",
X"18",
X"18",
X"3c",
X"00",
X"00",
X"00",
X"66",
X"7f",
X"7f",
X"6b",
X"63",
X"00",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"66",
X"66",
X"00",
X"00",
X"00",
X"3c",
X"66",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"7c",
X"60",
X"60",
X"00",
X"00",
X"3e",
X"66",
X"66",
X"3e",
X"06",
X"06",
X"00",
X"00",
X"7c",
X"66",
X"60",
X"60",
X"60",
X"00",
X"00",
X"00",
X"3e",
X"60",
X"3c",
X"06",
X"7c",
X"00",
X"00",
X"18",
X"7e",
X"18",
X"18",
X"18",
X"0e",
X"00",
X"00",
X"00",
X"66",
X"66",
X"66",
X"66",
X"3e",
X"00",
X"00",
X"00",
X"66",
X"66",
X"66",
X"3c",
X"18",
X"00",
X"00",
X"00",
X"63",
X"6b",
X"7f",
X"3e",
X"36",
X"00",
X"00",
X"00",
X"66",
X"3c",
X"18",
X"3c",
X"66",
X"00",
X"00",
X"00",
X"66",
X"66",
X"66",
X"3e",
X"0c",
X"78",
X"00",
X"00",
X"7e",
X"0c",
X"18",
X"30",
X"7e",
X"00",
X"00",
X"18",
X"3c",
X"7e",
X"7e",
X"18",
X"3c",
X"00",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"00",
X"7e",
X"78",
X"7c",
X"6e",
X"66",
X"06",
X"00",
X"08",
X"18",
X"38",
X"78",
X"38",
X"18",
X"08",
X"00",
X"10",
X"18",
X"1c",
X"1e",
X"1c",
X"18",
X"10",
X"00",
X"fb",
X"f3",
X"33",
X"f6",
X"3d",
X"f6",
X"a3",
X"f6",
X"33",
X"f6",
X"3c",
X"f6",
X"4c",
X"e4",
X"f3",
X"00",
X"f5",
X"f3",
X"33",
X"f6",
X"92",
X"f5",
X"b6",
X"f5",
X"33",
X"f6",
X"fb",
X"fc",
X"4c",
X"e4",
X"f3",
X"00",
X"33",
X"f6",
X"33",
X"f6",
X"e1",
X"f6",
X"3c",
X"f6",
X"33",
X"f6",
X"3c",
X"f6",
X"4c",
X"e4",
X"f3",
X"00",
X"9e",
X"ee",
X"db",
X"ee",
X"9d",
X"ee",
X"a6",
X"ee",
X"80",
X"ee",
X"9d",
X"ee",
X"4c",
X"78",
X"ee",
X"00",
X"4b",
X"ef",
X"2a",
X"f0",
X"d5",
X"ef",
X"0f",
X"f0",
X"27",
X"f0",
X"4a",
X"ef",
X"4c",
X"41",
X"ef",
X"00",
X"4c",
X"ea",
X"ed",
X"4c",
X"f0",
X"ed",
X"4c",
X"c4",
X"e4",
X"4c",
X"59",
X"e9",
X"4c",
X"ed",
X"e8",
X"4c",
X"ae",
X"e7",
X"4c",
X"05",
X"e9",
X"4c",
X"44",
X"e9",
X"4c",
X"f2",
X"eb",
X"4c",
X"d5",
X"e6",
X"4c",
X"a6",
X"e4",
X"4c",
X"23",
X"f2",
X"4c",
X"1b",
X"f1",
X"4c",
X"25",
X"f1",
X"4c",
X"e9",
X"ef",
X"4c",
X"5d",
X"ef",
X"90",
X"e7",
X"8f",
X"e7",
X"8f",
X"e7",
X"8f",
X"e7",
X"be",
X"ff",
X"0f",
X"eb",
X"90",
X"ea",
X"cf",
X"ea",
X"8f",
X"e7",
X"8f",
X"e7",
X"8f",
X"e7",
X"06",
X"e7",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ae",
X"e7",
X"05",
X"e9",
X"a2",
X"00",
X"a9",
X"ff",
X"9d",
X"40",
X"03",
X"a9",
X"c0",
X"9d",
X"46",
X"03",
X"a9",
X"e4",
X"9d",
X"47",
X"03",
X"8a",
X"18",
X"69",
X"10",
X"aa",
X"c9",
X"80",
X"90",
X"e8",
X"60",
X"a0",
X"85",
X"60",
X"85",
X"2f",
X"86",
X"2e",
X"8a",
X"29",
X"0f",
X"d0",
X"04",
X"e0",
X"80",
X"90",
X"05",
X"a0",
X"86",
X"4c",
X"1b",
X"e6",
X"a0",
X"00",
X"bd",
X"40",
X"03",
X"99",
X"20",
X"00",
X"e8",
X"c8",
X"c0",
X"0c",
X"90",
X"f4",
X"a0",
X"84",
X"a5",
X"22",
X"c9",
X"03",
X"90",
X"25",
X"a8",
X"c0",
X"0e",
X"90",
X"02",
X"a0",
X"0e",
X"84",
X"17",
X"b9",
X"c6",
X"e6",
X"f0",
X"0f",
X"c9",
X"02",
X"f0",
X"35",
X"c9",
X"08",
X"b0",
X"4c",
X"c9",
X"04",
X"f0",
X"63",
X"4c",
X"c9",
X"e5",
X"a5",
X"20",
X"c9",
X"ff",
X"f0",
X"05",
X"a0",
X"81",
X"4c",
X"1b",
X"e6",
X"20",
X"9e",
X"e6",
X"b0",
X"f8",
X"20",
X"3d",
X"e6",
X"b0",
X"f3",
X"20",
X"89",
X"e6",
X"a9",
X"0b",
X"85",
X"17",
X"20",
X"3d",
X"e6",
X"a5",
X"2c",
X"85",
X"26",
X"a5",
X"2d",
X"85",
X"27",
X"4c",
X"1d",
X"e6",
X"a0",
X"01",
X"84",
X"23",
X"20",
X"3d",
X"e6",
X"b0",
X"03",
X"20",
X"89",
X"e6",
X"a9",
X"ff",
X"85",
X"20",
X"a9",
X"e4",
X"85",
X"27",
X"a9",
X"c0",
X"85",
X"26",
X"4c",
X"1d",
X"e6",
X"a5",
X"20",
X"c9",
X"ff",
X"d0",
X"05",
X"20",
X"9e",
X"e6",
X"b0",
X"b8",
X"20",
X"3d",
X"e6",
X"20",
X"89",
X"e6",
X"a6",
X"2e",
X"bd",
X"40",
X"03",
X"85",
X"20",
X"4c",
X"1d",
X"e6",
X"a5",
X"22",
X"25",
X"2a",
X"d0",
X"05",
X"a0",
X"83",
X"4c",
X"1b",
X"e6",
X"20",
X"3d",
X"e6",
X"b0",
X"f8",
X"a5",
X"28",
X"05",
X"29",
X"d0",
X"08",
X"20",
X"89",
X"e6",
X"85",
X"2f",
X"4c",
X"1d",
X"e6",
X"20",
X"89",
X"e6",
X"85",
X"2f",
X"30",
X"35",
X"a0",
X"00",
X"91",
X"24",
X"20",
X"70",
X"e6",
X"a5",
X"22",
X"29",
X"02",
X"d0",
X"0c",
X"a5",
X"2f",
X"c9",
X"9b",
X"d0",
X"06",
X"20",
X"63",
X"e6",
X"4c",
X"c3",
X"e5",
X"20",
X"63",
X"e6",
X"d0",
X"db",
X"a5",
X"22",
X"29",
X"02",
X"d0",
X"11",
X"20",
X"89",
X"e6",
X"85",
X"2f",
X"30",
X"0a",
X"a5",
X"2f",
X"c9",
X"9b",
X"d0",
X"f3",
X"a9",
X"89",
X"85",
X"23",
X"20",
X"77",
X"e6",
X"4c",
X"1d",
X"e6",
X"a5",
X"22",
X"25",
X"2a",
X"d0",
X"05",
X"a0",
X"87",
X"4c",
X"1b",
X"e6",
X"20",
X"3d",
X"e6",
X"b0",
X"f8",
X"a5",
X"28",
X"05",
X"29",
X"d0",
X"06",
X"a5",
X"2f",
X"e6",
X"28",
X"d0",
X"06",
X"a0",
X"00",
X"b1",
X"24",
X"85",
X"2f",
X"20",
X"89",
X"e6",
X"30",
X"25",
X"20",
X"70",
X"e6",
X"a5",
X"22",
X"29",
X"02",
X"d0",
X"0c",
X"a5",
X"2f",
X"c9",
X"9b",
X"d0",
X"06",
X"20",
X"63",
X"e6",
X"4c",
X"15",
X"e6",
X"20",
X"63",
X"e6",
X"d0",
X"db",
X"a5",
X"22",
X"29",
X"02",
X"d0",
X"05",
X"a9",
X"9b",
X"20",
X"89",
X"e6",
X"20",
X"77",
X"e6",
X"4c",
X"1d",
X"e6",
X"84",
X"23",
X"a4",
X"2e",
X"b9",
X"44",
X"03",
X"85",
X"24",
X"b9",
X"45",
X"03",
X"85",
X"25",
X"a2",
X"00",
X"b5",
X"20",
X"99",
X"40",
X"03",
X"e8",
X"c8",
X"e0",
X"0c",
X"90",
X"f5",
X"a5",
X"2f",
X"a6",
X"2e",
X"a4",
X"23",
X"60",
X"a4",
X"20",
X"c0",
X"22",
X"90",
X"04",
X"a0",
X"85",
X"b0",
X"1b",
X"b9",
X"1b",
X"03",
X"85",
X"2c",
X"b9",
X"1c",
X"03",
X"85",
X"2d",
X"a4",
X"17",
X"b9",
X"c6",
X"e6",
X"a8",
X"b1",
X"2c",
X"aa",
X"c8",
X"b1",
X"2c",
X"85",
X"2d",
X"86",
X"2c",
X"18",
X"60",
X"c6",
X"28",
X"a5",
X"28",
X"c9",
X"ff",
X"d0",
X"02",
X"c6",
X"29",
X"05",
X"29",
X"60",
X"e6",
X"24",
X"d0",
X"02",
X"e6",
X"25",
X"60",
X"a6",
X"2e",
X"38",
X"bd",
X"48",
X"03",
X"e5",
X"28",
X"85",
X"28",
X"bd",
X"49",
X"03",
X"e5",
X"29",
X"85",
X"29",
X"60",
X"a0",
X"92",
X"20",
X"93",
X"e6",
X"84",
X"23",
X"c0",
X"00",
X"60",
X"aa",
X"a5",
X"2d",
X"48",
X"a5",
X"2c",
X"48",
X"8a",
X"a6",
X"2e",
X"60",
X"a0",
X"00",
X"b1",
X"24",
X"f0",
X"0c",
X"a0",
X"21",
X"d9",
X"1a",
X"03",
X"f0",
X"0a",
X"88",
X"88",
X"88",
X"10",
X"f6",
X"a0",
X"82",
X"38",
X"b0",
X"13",
X"98",
X"85",
X"20",
X"38",
X"a0",
X"01",
X"b1",
X"24",
X"e9",
X"30",
X"c9",
X"0a",
X"90",
X"02",
X"a9",
X"01",
X"85",
X"21",
X"18",
X"60",
X"00",
X"04",
X"04",
X"04",
X"04",
X"06",
X"06",
X"06",
X"06",
X"02",
X"08",
X"0a",
X"a9",
X"40",
X"8d",
X"0e",
X"d4",
X"a9",
X"38",
X"8d",
X"02",
X"d3",
X"8d",
X"03",
X"d3",
X"a9",
X"00",
X"8d",
X"00",
X"d3",
X"ea",
X"ea",
X"ea",
X"a9",
X"3c",
X"8d",
X"02",
X"d3",
X"8d",
X"03",
X"d3",
X"60",
X"6c",
X"16",
X"02",
X"80",
X"40",
X"04",
X"02",
X"01",
X"08",
X"10",
X"20",
X"36",
X"08",
X"14",
X"12",
X"10",
X"0e",
X"0c",
X"0a",
X"48",
X"ad",
X"0e",
X"d2",
X"29",
X"20",
X"d0",
X"0d",
X"a9",
X"df",
X"8d",
X"0e",
X"d2",
X"a5",
X"10",
X"8d",
X"0e",
X"d2",
X"6c",
X"0a",
X"02",
X"8a",
X"48",
X"a2",
X"06",
X"bd",
X"f6",
X"e6",
X"e0",
X"05",
X"d0",
X"04",
X"25",
X"10",
X"f0",
X"05",
X"2c",
X"0e",
X"d2",
X"f0",
X"06",
X"ca",
X"10",
X"ed",
X"4c",
X"62",
X"e7",
X"49",
X"ff",
X"8d",
X"0e",
X"d2",
X"a5",
X"10",
X"8d",
X"0e",
X"d2",
X"bd",
X"fe",
X"e6",
X"aa",
X"bd",
X"00",
X"02",
X"8d",
X"8c",
X"02",
X"bd",
X"01",
X"02",
X"8d",
X"8d",
X"02",
X"68",
X"aa",
X"6c",
X"8c",
X"02",
X"a9",
X"00",
X"85",
X"11",
X"8d",
X"ff",
X"02",
X"8d",
X"f0",
X"02",
X"85",
X"4d",
X"68",
X"40",
X"68",
X"aa",
X"2c",
X"02",
X"d3",
X"10",
X"06",
X"ad",
X"00",
X"d3",
X"6c",
X"02",
X"02",
X"2c",
X"03",
X"d3",
X"10",
X"06",
X"ad",
X"01",
X"d3",
X"6c",
X"04",
X"02",
X"68",
X"8d",
X"8c",
X"02",
X"68",
X"48",
X"29",
X"10",
X"f0",
X"07",
X"ad",
X"8c",
X"02",
X"48",
X"6c",
X"06",
X"02",
X"ad",
X"8c",
X"02",
X"48",
X"68",
X"40",
X"2c",
X"0f",
X"d4",
X"10",
X"03",
X"6c",
X"00",
X"02",
X"48",
X"ad",
X"0f",
X"d4",
X"29",
X"20",
X"f0",
X"03",
X"4c",
X"74",
X"e4",
X"8a",
X"48",
X"98",
X"48",
X"8d",
X"0f",
X"d4",
X"6c",
X"22",
X"02",
X"e6",
X"14",
X"d0",
X"08",
X"e6",
X"4d",
X"e6",
X"13",
X"d0",
X"02",
X"e6",
X"12",
X"a9",
X"fe",
X"a2",
X"00",
X"a4",
X"4d",
X"10",
X"06",
X"85",
X"4d",
X"a6",
X"13",
X"a9",
X"f6",
X"85",
X"4e",
X"86",
X"4f",
X"a2",
X"00",
X"20",
X"d0",
X"e8",
X"d0",
X"03",
X"20",
X"ca",
X"e8",
X"a5",
X"42",
X"d0",
X"08",
X"ba",
X"bd",
X"04",
X"01",
X"29",
X"04",
X"f0",
X"03",
X"4c",
X"05",
X"e9",
X"ad",
X"0d",
X"d4",
X"8d",
X"35",
X"02",
X"ad",
X"0c",
X"d4",
X"8d",
X"34",
X"02",
X"ad",
X"31",
X"02",
X"8d",
X"03",
X"d4",
X"ad",
X"30",
X"02",
X"8d",
X"02",
X"d4",
X"ad",
X"2f",
X"02",
X"8d",
X"00",
X"d4",
X"ad",
X"6f",
X"02",
X"8d",
X"1b",
X"d0",
X"a2",
X"08",
X"8e",
X"1f",
X"d0",
X"58",
X"bd",
X"c0",
X"02",
X"45",
X"4f",
X"25",
X"4e",
X"9d",
X"12",
X"d0",
X"ca",
X"10",
X"f2",
X"ad",
X"f4",
X"02",
X"8d",
X"09",
X"d4",
X"ad",
X"f3",
X"02",
X"8d",
X"01",
X"d4",
X"a2",
X"02",
X"20",
X"d0",
X"e8",
X"d0",
X"03",
X"20",
X"cd",
X"e8",
X"a2",
X"02",
X"e8",
X"e8",
X"bd",
X"18",
X"02",
X"1d",
X"19",
X"02",
X"f0",
X"06",
X"20",
X"d0",
X"e8",
X"9d",
X"26",
X"02",
X"e0",
X"08",
X"d0",
X"ec",
X"ad",
X"0f",
X"d2",
X"29",
X"04",
X"f0",
X"08",
X"ad",
X"f1",
X"02",
X"f0",
X"03",
X"ce",
X"f1",
X"02",
X"ad",
X"2b",
X"02",
X"f0",
X"17",
X"ad",
X"0f",
X"d2",
X"29",
X"04",
X"d0",
X"60",
X"ce",
X"2b",
X"02",
X"d0",
X"0b",
X"a9",
X"06",
X"8d",
X"2b",
X"02",
X"ad",
X"09",
X"d2",
X"8d",
X"fc",
X"02",
X"a0",
X"01",
X"a2",
X"03",
X"b9",
X"00",
X"d3",
X"4a",
X"4a",
X"4a",
X"4a",
X"9d",
X"78",
X"02",
X"ca",
X"b9",
X"00",
X"d3",
X"29",
X"0f",
X"9d",
X"78",
X"02",
X"ca",
X"88",
X"10",
X"e9",
X"a2",
X"03",
X"bd",
X"10",
X"d0",
X"9d",
X"84",
X"02",
X"bd",
X"00",
X"d2",
X"9d",
X"70",
X"02",
X"bd",
X"04",
X"d2",
X"9d",
X"74",
X"02",
X"ca",
X"10",
X"eb",
X"8d",
X"0b",
X"d2",
X"a2",
X"06",
X"a0",
X"03",
X"b9",
X"78",
X"02",
X"4a",
X"4a",
X"4a",
X"9d",
X"7d",
X"02",
X"a9",
X"00",
X"2a",
X"9d",
X"7c",
X"02",
X"ca",
X"ca",
X"88",
X"10",
X"ec",
X"6c",
X"24",
X"02",
X"a9",
X"00",
X"8d",
X"2b",
X"02",
X"f0",
X"a9",
X"6c",
X"26",
X"02",
X"6c",
X"28",
X"02",
X"bc",
X"18",
X"02",
X"d0",
X"08",
X"bc",
X"19",
X"02",
X"f0",
X"10",
X"de",
X"19",
X"02",
X"de",
X"18",
X"02",
X"d0",
X"08",
X"bc",
X"19",
X"02",
X"d0",
X"03",
X"a9",
X"00",
X"60",
X"a9",
X"ff",
X"60",
X"0a",
X"8d",
X"2d",
X"02",
X"8a",
X"a2",
X"05",
X"8d",
X"0a",
X"d4",
X"ca",
X"d0",
X"fd",
X"ae",
X"2d",
X"02",
X"9d",
X"17",
X"02",
X"98",
X"9d",
X"16",
X"02",
X"60",
X"68",
X"a8",
X"68",
X"aa",
X"68",
X"40",
X"66",
X"66",
X"7e",
X"66",
X"00",
X"00",
X"7c",
X"4c",
X"ed",
X"e8",
X"66",
X"7c",
X"00",
X"00",
X"3c",
X"66",
X"60",
X"60",
X"66",
X"3c",
X"00",
X"00",
X"78",
X"6c",
X"66",
X"66",
X"6c",
X"78",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"60",
X"60",
X"7e",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"60",
X"60",
X"60",
X"00",
X"00",
X"3e",
X"60",
X"60",
X"6e",
X"66",
X"3e",
X"00",
X"00",
X"66",
X"66",
X"7e",
X"a9",
X"3c",
X"8d",
X"02",
X"d3",
X"a9",
X"3c",
X"8d",
X"03",
X"d3",
X"a9",
X"03",
X"8d",
X"32",
X"02",
X"85",
X"41",
X"8d",
X"0f",
X"d2",
X"60",
X"ba",
X"8e",
X"18",
X"03",
X"a9",
X"01",
X"85",
X"42",
X"ad",
X"00",
X"03",
X"c9",
X"60",
X"d0",
X"03",
X"4c",
X"80",
X"eb",
X"a9",
X"00",
X"8d",
X"0f",
X"03",
X"a9",
X"01",
X"85",
X"37",
X"a9",
X"0d",
X"85",
X"36",
X"a9",
X"28",
X"8d",
X"04",
X"d2",
X"a9",
X"00",
X"8d",
X"06",
X"d2",
X"18",
X"ad",
X"00",
X"03",
X"6d",
X"01",
X"03",
X"69",
X"ff",
X"8d",
X"3a",
X"02",
X"ad",
X"02",
X"03",
X"8d",
X"3b",
X"02",
X"ad",
X"0a",
X"03",
X"8d",
X"3c",
X"02",
X"ad",
X"0b",
X"03",
X"8d",
X"3d",
X"02",
X"18",
X"a9",
X"3a",
X"85",
X"32",
X"69",
X"04",
X"85",
X"34",
X"a9",
X"02",
X"85",
X"33",
X"85",
X"35",
X"a9",
X"34",
X"8d",
X"03",
X"d3",
X"20",
X"8a",
X"ec",
X"ad",
X"3f",
X"02",
X"d0",
X"03",
X"98",
X"d0",
X"07",
X"c6",
X"36",
X"10",
X"b5",
X"4c",
X"06",
X"ea",
X"ad",
X"03",
X"03",
X"10",
X"0c",
X"a9",
X"0d",
X"85",
X"36",
X"20",
X"6a",
X"eb",
X"20",
X"8a",
X"ec",
X"f0",
X"e8",
X"20",
X"75",
X"ec",
X"a9",
X"00",
X"8d",
X"3f",
X"02",
X"20",
X"9b",
X"ec",
X"f0",
X"12",
X"2c",
X"03",
X"03",
X"70",
X"07",
X"ad",
X"3f",
X"02",
X"d0",
X"18",
X"f0",
X"1d",
X"20",
X"6a",
X"eb",
X"20",
X"e0",
X"ea",
X"ad",
X"3f",
X"02",
X"f0",
X"05",
X"ad",
X"19",
X"03",
X"85",
X"30",
X"a5",
X"30",
X"c9",
X"01",
X"f0",
X"07",
X"c6",
X"37",
X"30",
X"03",
X"4c",
X"74",
X"e9",
X"20",
X"5f",
X"ec",
X"a9",
X"00",
X"85",
X"42",
X"a4",
X"30",
X"8c",
X"03",
X"03",
X"60",
X"a9",
X"00",
X"8d",
X"3f",
X"02",
X"18",
X"a9",
X"3e",
X"85",
X"32",
X"69",
X"01",
X"85",
X"34",
X"a9",
X"02",
X"85",
X"33",
X"85",
X"35",
X"a9",
X"ff",
X"85",
X"3c",
X"20",
X"e0",
X"ea",
X"a0",
X"ff",
X"a5",
X"30",
X"c9",
X"01",
X"d0",
X"19",
X"ad",
X"3e",
X"02",
X"c9",
X"41",
X"f0",
X"21",
X"c9",
X"43",
X"f0",
X"1d",
X"c9",
X"45",
X"d0",
X"06",
X"a9",
X"90",
X"85",
X"30",
X"d0",
X"04",
X"a9",
X"8b",
X"85",
X"30",
X"a5",
X"30",
X"c9",
X"8a",
X"f0",
X"07",
X"a9",
X"ff",
X"8d",
X"3f",
X"02",
X"d0",
X"02",
X"a0",
X"00",
X"a5",
X"30",
X"8d",
X"19",
X"03",
X"60",
X"a9",
X"01",
X"85",
X"30",
X"20",
X"f2",
X"eb",
X"a0",
X"00",
X"84",
X"31",
X"84",
X"3b",
X"84",
X"3a",
X"b1",
X"32",
X"8d",
X"0d",
X"d2",
X"85",
X"31",
X"a5",
X"11",
X"d0",
X"03",
X"4c",
X"a0",
X"ed",
X"a5",
X"3a",
X"f0",
X"f5",
X"20",
X"5f",
X"ec",
X"60",
X"98",
X"48",
X"e6",
X"32",
X"d0",
X"02",
X"e6",
X"33",
X"a5",
X"32",
X"c5",
X"34",
X"a5",
X"33",
X"e5",
X"35",
X"90",
X"1c",
X"a5",
X"3b",
X"d0",
X"0b",
X"a5",
X"31",
X"8d",
X"0d",
X"d2",
X"a9",
X"ff",
X"85",
X"3b",
X"d0",
X"09",
X"a5",
X"10",
X"09",
X"08",
X"85",
X"10",
X"8d",
X"0e",
X"d2",
X"68",
X"a8",
X"68",
X"40",
X"a0",
X"00",
X"b1",
X"32",
X"8d",
X"0d",
X"d2",
X"18",
X"65",
X"31",
X"69",
X"00",
X"85",
X"31",
X"4c",
X"ba",
X"ea",
X"a5",
X"3b",
X"f0",
X"0b",
X"85",
X"3a",
X"a5",
X"10",
X"29",
X"f7",
X"85",
X"10",
X"8d",
X"0e",
X"d2",
X"68",
X"40",
X"a9",
X"00",
X"ac",
X"0f",
X"03",
X"d0",
X"02",
X"85",
X"31",
X"85",
X"38",
X"85",
X"39",
X"a9",
X"01",
X"85",
X"30",
X"20",
X"1b",
X"ec",
X"a9",
X"3c",
X"8d",
X"03",
X"d3",
X"a5",
X"11",
X"d0",
X"03",
X"4c",
X"a0",
X"ed",
X"ad",
X"17",
X"03",
X"f0",
X"05",
X"a5",
X"39",
X"f0",
X"f0",
X"60",
X"a9",
X"8a",
X"85",
X"30",
X"60",
X"98",
X"48",
X"ad",
X"0f",
X"d2",
X"8d",
X"0a",
X"d2",
X"30",
X"04",
X"a0",
X"8c",
X"84",
X"30",
X"29",
X"20",
X"d0",
X"04",
X"a0",
X"8e",
X"84",
X"30",
X"a5",
X"38",
X"f0",
X"13",
X"ad",
X"0d",
X"d2",
X"c5",
X"31",
X"f0",
X"04",
X"a0",
X"8f",
X"84",
X"30",
X"a9",
X"ff",
X"85",
X"39",
X"68",
X"a8",
X"68",
X"40",
X"ad",
X"0d",
X"d2",
X"a0",
X"00",
X"91",
X"32",
X"18",
X"65",
X"31",
X"69",
X"00",
X"85",
X"31",
X"e6",
X"32",
X"d0",
X"02",
X"e6",
X"33",
X"a5",
X"32",
X"c5",
X"34",
X"a5",
X"33",
X"e5",
X"35",
X"90",
X"de",
X"a5",
X"3c",
X"f0",
X"06",
X"a9",
X"00",
X"85",
X"3c",
X"f0",
X"d0",
X"a9",
X"ff",
X"85",
X"38",
X"d0",
X"ce",
X"18",
X"ad",
X"04",
X"03",
X"85",
X"32",
X"6d",
X"08",
X"03",
X"85",
X"34",
X"ad",
X"05",
X"03",
X"85",
X"33",
X"6d",
X"09",
X"03",
X"85",
X"35",
X"60",
X"ad",
X"03",
X"03",
X"10",
X"2e",
X"a9",
X"cc",
X"8d",
X"04",
X"d2",
X"a9",
X"05",
X"8d",
X"06",
X"d2",
X"20",
X"f2",
X"eb",
X"a0",
X"0f",
X"ad",
X"0b",
X"03",
X"30",
X"02",
X"a0",
X"b4",
X"a2",
X"00",
X"20",
X"b9",
X"ed",
X"a9",
X"34",
X"8d",
X"02",
X"d3",
X"ad",
X"17",
X"03",
X"d0",
X"fb",
X"20",
X"6a",
X"eb",
X"20",
X"6b",
X"ea",
X"4c",
X"df",
X"eb",
X"a9",
X"ff",
X"8d",
X"0f",
X"03",
X"a0",
X"0a",
X"ad",
X"0b",
X"03",
X"30",
X"02",
X"a0",
X"78",
X"a2",
X"00",
X"20",
X"b9",
X"ed",
X"a9",
X"34",
X"8d",
X"02",
X"d3",
X"ad",
X"17",
X"03",
X"d0",
X"fb",
X"20",
X"6a",
X"eb",
X"20",
X"75",
X"ec",
X"20",
X"b9",
X"ed",
X"20",
X"10",
X"ed",
X"20",
X"e0",
X"ea",
X"ad",
X"0b",
X"03",
X"30",
X"05",
X"a9",
X"3c",
X"8d",
X"02",
X"d3",
X"4c",
X"0d",
X"ea",
X"a9",
X"00",
X"8d",
X"17",
X"03",
X"60",
X"a9",
X"07",
X"2d",
X"32",
X"02",
X"09",
X"20",
X"ac",
X"00",
X"03",
X"c0",
X"60",
X"d0",
X"0c",
X"09",
X"08",
X"a0",
X"07",
X"8c",
X"02",
X"d2",
X"a0",
X"05",
X"8c",
X"00",
X"d2",
X"8d",
X"32",
X"02",
X"8d",
X"0f",
X"d2",
X"a9",
X"c7",
X"25",
X"10",
X"09",
X"10",
X"4c",
X"31",
X"ec",
X"a9",
X"07",
X"2d",
X"32",
X"02",
X"09",
X"10",
X"8d",
X"32",
X"02",
X"8d",
X"0f",
X"d2",
X"8d",
X"0a",
X"d2",
X"a9",
X"c7",
X"25",
X"10",
X"09",
X"20",
X"85",
X"10",
X"8d",
X"0e",
X"d2",
X"a9",
X"28",
X"8d",
X"08",
X"d2",
X"a2",
X"06",
X"a9",
X"a8",
X"a4",
X"41",
X"d0",
X"02",
X"a9",
X"a0",
X"9d",
X"01",
X"d2",
X"ca",
X"ca",
X"10",
X"f9",
X"a9",
X"a0",
X"8d",
X"05",
X"d2",
X"ac",
X"00",
X"03",
X"c0",
X"60",
X"f0",
X"06",
X"8d",
X"01",
X"d2",
X"8d",
X"03",
X"d2",
X"60",
X"ea",
X"a9",
X"c7",
X"25",
X"10",
X"85",
X"10",
X"8d",
X"0e",
X"d2",
X"a2",
X"06",
X"a9",
X"00",
X"9d",
X"01",
X"d2",
X"ca",
X"ca",
X"10",
X"f9",
X"60",
X"ad",
X"06",
X"03",
X"6a",
X"6a",
X"a8",
X"29",
X"3f",
X"aa",
X"98",
X"6a",
X"29",
X"c0",
X"a8",
X"60",
X"0f",
X"eb",
X"90",
X"ea",
X"cf",
X"ea",
X"a2",
X"01",
X"a0",
X"ff",
X"88",
X"d0",
X"fd",
X"ca",
X"d0",
X"f8",
X"20",
X"6b",
X"ea",
X"a0",
X"02",
X"a2",
X"00",
X"20",
X"b9",
X"ed",
X"20",
X"1a",
X"ea",
X"98",
X"60",
X"8d",
X"10",
X"03",
X"8c",
X"11",
X"03",
X"20",
X"04",
X"ed",
X"8d",
X"10",
X"03",
X"ad",
X"0c",
X"03",
X"20",
X"04",
X"ed",
X"8d",
X"0c",
X"03",
X"ad",
X"10",
X"03",
X"38",
X"ed",
X"0c",
X"03",
X"8d",
X"12",
X"03",
X"ad",
X"11",
X"03",
X"38",
X"ed",
X"0d",
X"03",
X"a8",
X"a9",
X"7d",
X"18",
X"69",
X"83",
X"88",
X"10",
X"fa",
X"18",
X"6d",
X"12",
X"03",
X"a8",
X"4a",
X"4a",
X"4a",
X"0a",
X"38",
X"e9",
X"16",
X"aa",
X"98",
X"29",
X"07",
X"a8",
X"a9",
X"f5",
X"18",
X"69",
X"0b",
X"88",
X"10",
X"fa",
X"a0",
X"00",
X"8c",
X"0e",
X"03",
X"38",
X"e9",
X"07",
X"10",
X"03",
X"ce",
X"0e",
X"03",
X"18",
X"7d",
X"d0",
X"ed",
X"a8",
X"ad",
X"0e",
X"03",
X"7d",
X"d1",
X"ed",
X"60",
X"c9",
X"7c",
X"30",
X"04",
X"38",
X"e9",
X"7c",
X"60",
X"18",
X"69",
X"07",
X"60",
X"a5",
X"11",
X"d0",
X"03",
X"4c",
X"a0",
X"ed",
X"78",
X"ad",
X"17",
X"03",
X"d0",
X"02",
X"f0",
X"25",
X"ad",
X"0f",
X"d2",
X"29",
X"10",
X"d0",
X"ea",
X"8d",
X"16",
X"03",
X"ae",
X"0b",
X"d4",
X"a4",
X"14",
X"8e",
X"0c",
X"03",
X"8c",
X"0d",
X"03",
X"a2",
X"01",
X"8e",
X"15",
X"03",
X"a0",
X"0a",
X"a5",
X"11",
X"f0",
X"61",
X"ad",
X"17",
X"03",
X"d0",
X"04",
X"58",
X"4c",
X"0a",
X"eb",
X"ad",
X"0f",
X"d2",
X"29",
X"10",
X"cd",
X"16",
X"03",
X"f0",
X"e9",
X"8d",
X"16",
X"03",
X"88",
X"d0",
X"e3",
X"ce",
X"15",
X"03",
X"30",
X"12",
X"ad",
X"0b",
X"d4",
X"a4",
X"14",
X"20",
X"a3",
X"ec",
X"8c",
X"ee",
X"02",
X"8d",
X"ef",
X"02",
X"a0",
X"09",
X"d0",
X"cc",
X"ad",
X"ee",
X"02",
X"8d",
X"04",
X"d2",
X"ad",
X"ef",
X"02",
X"8d",
X"06",
X"d2",
X"a9",
X"00",
X"8d",
X"0f",
X"d2",
X"ad",
X"32",
X"02",
X"8d",
X"0f",
X"d2",
X"a9",
X"55",
X"91",
X"32",
X"c8",
X"91",
X"32",
X"a9",
X"aa",
X"85",
X"31",
X"18",
X"a5",
X"32",
X"69",
X"02",
X"85",
X"32",
X"a5",
X"33",
X"69",
X"00",
X"85",
X"33",
X"58",
X"60",
X"20",
X"5f",
X"ec",
X"a9",
X"3c",
X"8d",
X"02",
X"d3",
X"8d",
X"03",
X"d3",
X"a9",
X"80",
X"85",
X"30",
X"ae",
X"18",
X"03",
X"9a",
X"c6",
X"11",
X"58",
X"4c",
X"0d",
X"ea",
X"a9",
X"ec",
X"8d",
X"26",
X"02",
X"a9",
X"eb",
X"8d",
X"27",
X"02",
X"a9",
X"01",
X"78",
X"20",
X"5c",
X"e4",
X"a9",
X"01",
X"8d",
X"17",
X"03",
X"58",
X"60",
X"e8",
X"03",
X"43",
X"04",
X"9e",
X"04",
X"f9",
X"04",
X"54",
X"05",
X"af",
X"05",
X"0a",
X"06",
X"65",
X"06",
X"c0",
X"06",
X"1a",
X"07",
X"75",
X"07",
X"d0",
X"07",
X"24",
X"85",
X"a9",
X"a0",
X"8d",
X"46",
X"02",
X"60",
X"a9",
X"31",
X"8d",
X"00",
X"03",
X"ad",
X"46",
X"02",
X"ae",
X"02",
X"03",
X"e0",
X"21",
X"f0",
X"02",
X"a9",
X"07",
X"8d",
X"06",
X"03",
X"a2",
X"40",
X"a0",
X"80",
X"ad",
X"02",
X"03",
X"c9",
X"57",
X"d0",
X"02",
X"a2",
X"80",
X"c9",
X"53",
X"d0",
X"0c",
X"a9",
X"ea",
X"8d",
X"04",
X"03",
X"a9",
X"02",
X"8d",
X"05",
X"03",
X"a0",
X"04",
X"8e",
X"03",
X"03",
X"8c",
X"08",
X"03",
X"a9",
X"00",
X"8d",
X"09",
X"03",
X"20",
X"59",
X"e4",
X"10",
X"01",
X"60",
X"ad",
X"02",
X"03",
X"c9",
X"53",
X"d0",
X"0a",
X"20",
X"6d",
X"ee",
X"a0",
X"02",
X"b1",
X"15",
X"8d",
X"46",
X"02",
X"ad",
X"02",
X"03",
X"c9",
X"21",
X"d0",
X"1f",
X"20",
X"6d",
X"ee",
X"a0",
X"fe",
X"c8",
X"c8",
X"b1",
X"15",
X"c9",
X"ff",
X"d0",
X"f8",
X"c8",
X"b1",
X"15",
X"c8",
X"c9",
X"ff",
X"d0",
X"f2",
X"88",
X"88",
X"8c",
X"08",
X"03",
X"a9",
X"00",
X"8d",
X"09",
X"03",
X"ac",
X"03",
X"03",
X"60",
X"ad",
X"04",
X"03",
X"85",
X"15",
X"ad",
X"05",
X"03",
X"85",
X"16",
X"60",
X"a9",
X"1e",
X"85",
X"1c",
X"60",
X"ea",
X"02",
X"c0",
X"03",
X"a9",
X"04",
X"85",
X"1e",
X"ae",
X"7d",
X"ee",
X"ac",
X"7e",
X"ee",
X"a9",
X"53",
X"8d",
X"02",
X"03",
X"8d",
X"0a",
X"03",
X"20",
X"e6",
X"ee",
X"20",
X"59",
X"e4",
X"30",
X"03",
X"20",
X"14",
X"ef",
X"60",
X"20",
X"81",
X"ee",
X"a9",
X"00",
X"85",
X"1d",
X"60",
X"85",
X"1f",
X"20",
X"1a",
X"ef",
X"a6",
X"1d",
X"a5",
X"1f",
X"9d",
X"c0",
X"03",
X"e8",
X"e4",
X"1e",
X"f0",
X"13",
X"86",
X"1d",
X"c9",
X"9b",
X"f0",
X"03",
X"a0",
X"01",
X"60",
X"a9",
X"20",
X"9d",
X"c0",
X"03",
X"e8",
X"e4",
X"1e",
X"d0",
X"f8",
X"a9",
X"00",
X"85",
X"1d",
X"ae",
X"7f",
X"ee",
X"ac",
X"80",
X"ee",
X"20",
X"e6",
X"ee",
X"20",
X"59",
X"e4",
X"60",
X"20",
X"1a",
X"ef",
X"a6",
X"1d",
X"d0",
X"de",
X"a0",
X"01",
X"60",
X"8e",
X"04",
X"03",
X"8c",
X"05",
X"03",
X"a9",
X"40",
X"8d",
X"00",
X"03",
X"a9",
X"01",
X"8d",
X"01",
X"03",
X"a9",
X"80",
X"ae",
X"02",
X"03",
X"e0",
X"53",
X"d0",
X"02",
X"a9",
X"40",
X"8d",
X"03",
X"03",
X"a5",
X"1e",
X"8d",
X"08",
X"03",
X"a9",
X"00",
X"8d",
X"09",
X"03",
X"a5",
X"1c",
X"8d",
X"06",
X"03",
X"60",
X"ad",
X"ec",
X"02",
X"85",
X"1c",
X"60",
X"a0",
X"57",
X"a5",
X"2b",
X"c9",
X"4e",
X"d0",
X"04",
X"a2",
X"28",
X"d0",
X"0e",
X"c9",
X"44",
X"d0",
X"04",
X"a2",
X"14",
X"d0",
X"06",
X"c9",
X"53",
X"d0",
X"0b",
X"a2",
X"1d",
X"86",
X"1e",
X"8c",
X"02",
X"03",
X"8d",
X"0a",
X"03",
X"60",
X"a9",
X"4e",
X"d0",
X"dd",
X"a9",
X"cc",
X"8d",
X"ee",
X"02",
X"a9",
X"05",
X"8d",
X"ef",
X"02",
X"60",
X"a5",
X"2b",
X"85",
X"3e",
X"a5",
X"2a",
X"29",
X"0c",
X"c9",
X"04",
X"f0",
X"05",
X"c9",
X"08",
X"f0",
X"39",
X"60",
X"a9",
X"00",
X"8d",
X"89",
X"02",
X"85",
X"3f",
X"a9",
X"01",
X"20",
X"58",
X"f0",
X"30",
X"24",
X"a9",
X"34",
X"8d",
X"02",
X"d3",
X"a0",
X"40",
X"a2",
X"02",
X"a9",
X"03",
X"8d",
X"2a",
X"02",
X"20",
X"5c",
X"e4",
X"ad",
X"2a",
X"02",
X"d0",
X"fb",
X"a9",
X"80",
X"85",
X"3d",
X"8d",
X"8a",
X"02",
X"4c",
X"d3",
X"ef",
X"a0",
X"80",
X"c6",
X"11",
X"a9",
X"00",
X"8d",
X"89",
X"02",
X"60",
X"a9",
X"80",
X"8d",
X"89",
X"02",
X"a9",
X"02",
X"20",
X"58",
X"f0",
X"30",
X"ee",
X"a9",
X"cc",
X"8d",
X"04",
X"d2",
X"a9",
X"05",
X"8d",
X"06",
X"d2",
X"a9",
X"60",
X"8d",
X"00",
X"03",
X"20",
X"68",
X"e4",
X"a9",
X"34",
X"8d",
X"02",
X"d3",
X"a9",
X"03",
X"a2",
X"04",
X"a0",
X"80",
X"20",
X"5c",
X"e4",
X"a9",
X"ff",
X"8d",
X"2a",
X"02",
X"a5",
X"11",
X"f0",
X"c1",
X"ad",
X"2a",
X"02",
X"d0",
X"f7",
X"a9",
X"00",
X"85",
X"3d",
X"a0",
X"01",
X"60",
X"a5",
X"3f",
X"30",
X"33",
X"a6",
X"3d",
X"ec",
X"8a",
X"02",
X"f0",
X"08",
X"bd",
X"00",
X"04",
X"e6",
X"3d",
X"a0",
X"01",
X"60",
X"a9",
X"52",
X"20",
X"95",
X"f0",
X"98",
X"30",
X"f7",
X"a9",
X"00",
X"85",
X"3d",
X"a2",
X"80",
X"ad",
X"ff",
X"03",
X"c9",
X"fe",
X"f0",
X"0d",
X"c9",
X"fa",
X"d0",
X"03",
X"ae",
X"7f",
X"04",
X"8e",
X"8a",
X"02",
X"4c",
X"d6",
X"ef",
X"c6",
X"3f",
X"a0",
X"88",
X"60",
X"a6",
X"3d",
X"9d",
X"00",
X"04",
X"e6",
X"3d",
X"a0",
X"01",
X"e0",
X"7f",
X"f0",
X"01",
X"60",
X"a9",
X"fc",
X"20",
X"d2",
X"f0",
X"a9",
X"00",
X"85",
X"3d",
X"60",
X"a0",
X"01",
X"60",
X"ad",
X"89",
X"02",
X"30",
X"08",
X"a0",
X"01",
X"a9",
X"3c",
X"8d",
X"02",
X"d3",
X"60",
X"a6",
X"3d",
X"f0",
X"0a",
X"8e",
X"7f",
X"04",
X"a9",
X"fa",
X"20",
X"d2",
X"f0",
X"30",
X"ec",
X"a2",
X"7f",
X"a9",
X"00",
X"9d",
X"00",
X"04",
X"ca",
X"10",
X"fa",
X"a9",
X"fe",
X"20",
X"d2",
X"f0",
X"4c",
X"32",
X"f0",
X"85",
X"40",
X"a5",
X"14",
X"18",
X"69",
X"1e",
X"aa",
X"a9",
X"ff",
X"8d",
X"1f",
X"d0",
X"a9",
X"00",
X"a0",
X"f0",
X"88",
X"d0",
X"fd",
X"8d",
X"1f",
X"d0",
X"a0",
X"f0",
X"88",
X"d0",
X"fd",
X"e4",
X"14",
X"d0",
X"e8",
X"c6",
X"40",
X"f0",
X"0b",
X"8a",
X"18",
X"69",
X"0a",
X"aa",
X"e4",
X"14",
X"d0",
X"fc",
X"f0",
X"d3",
X"20",
X"8c",
X"f0",
X"98",
X"60",
X"ad",
X"25",
X"e4",
X"48",
X"ad",
X"24",
X"e4",
X"48",
X"60",
X"8d",
X"02",
X"03",
X"a9",
X"00",
X"8d",
X"09",
X"03",
X"a9",
X"83",
X"8d",
X"08",
X"03",
X"a9",
X"03",
X"8d",
X"05",
X"03",
X"a9",
X"fd",
X"8d",
X"04",
X"03",
X"a9",
X"60",
X"8d",
X"00",
X"03",
X"a9",
X"00",
X"8d",
X"01",
X"03",
X"a9",
X"23",
X"8d",
X"06",
X"03",
X"ad",
X"02",
X"03",
X"a0",
X"40",
X"c9",
X"52",
X"f0",
X"02",
X"a0",
X"80",
X"8c",
X"03",
X"03",
X"a5",
X"3e",
X"8d",
X"0b",
X"03",
X"20",
X"59",
X"e4",
X"60",
X"8d",
X"ff",
X"03",
X"a9",
X"55",
X"8d",
X"fd",
X"03",
X"8d",
X"fe",
X"03",
X"a9",
X"57",
X"20",
X"95",
X"f0",
X"60",
X"50",
X"30",
X"e4",
X"43",
X"40",
X"e4",
X"45",
X"00",
X"e4",
X"53",
X"10",
X"e4",
X"4b",
X"20",
X"e4",
X"7d",
X"41",
X"54",
X"41",
X"52",
X"49",
X"20",
X"43",
X"4f",
X"4d",
X"50",
X"55",
X"54",
X"45",
X"52",
X"20",
X"2d",
X"20",
X"4d",
X"45",
X"4d",
X"4f",
X"20",
X"50",
X"41",
X"44",
X"9b",
X"42",
X"4f",
X"4f",
X"54",
X"20",
X"45",
X"52",
X"52",
X"4f",
X"52",
X"9b",
X"45",
X"3a",
X"9b",
X"78",
X"ad",
X"44",
X"02",
X"d0",
X"04",
X"a9",
X"ff",
X"d0",
X"03",
X"78",
X"a9",
X"00",
X"85",
X"08",
X"d8",
X"a2",
X"ff",
X"9a",
X"20",
X"44",
X"f2",
X"20",
X"77",
X"f2",
X"a5",
X"08",
X"d0",
X"28",
X"a9",
X"00",
X"a0",
X"08",
X"85",
X"04",
X"85",
X"05",
X"91",
X"04",
X"c8",
X"c0",
X"00",
X"d0",
X"f9",
X"e6",
X"05",
X"a6",
X"05",
X"e4",
X"06",
X"d0",
X"f1",
X"ad",
X"72",
X"e4",
X"85",
X"0a",
X"ad",
X"73",
X"e4",
X"85",
X"0b",
X"a9",
X"ff",
X"8d",
X"44",
X"02",
X"d0",
X"13",
X"a2",
X"00",
X"8a",
X"9d",
X"00",
X"02",
X"9d",
X"00",
X"03",
X"ca",
X"d0",
X"f7",
X"a2",
X"10",
X"95",
X"00",
X"e8",
X"10",
X"fb",
X"a9",
X"02",
X"85",
X"52",
X"a9",
X"27",
X"85",
X"53",
X"a2",
X"25",
X"bd",
X"80",
X"e4",
X"9d",
X"00",
X"02",
X"ca",
X"10",
X"f7",
X"20",
X"8a",
X"f2",
X"58",
X"a2",
X"0e",
X"bd",
X"e3",
X"f0",
X"9d",
X"1a",
X"03",
X"ca",
X"10",
X"f7",
X"a2",
X"00",
X"86",
X"07",
X"86",
X"06",
X"ae",
X"e4",
X"02",
X"e0",
X"90",
X"b0",
X"0a",
X"ad",
X"fc",
X"9f",
X"d0",
X"05",
X"e6",
X"07",
X"20",
X"3c",
X"f2",
X"ae",
X"e4",
X"02",
X"e0",
X"b0",
X"b0",
X"0a",
X"ae",
X"fc",
X"bf",
X"d0",
X"05",
X"e6",
X"06",
X"20",
X"39",
X"f2",
X"a9",
X"03",
X"a2",
X"00",
X"9d",
X"42",
X"03",
X"a9",
X"18",
X"9d",
X"44",
X"03",
X"a9",
X"f1",
X"9d",
X"45",
X"03",
X"a9",
X"0c",
X"9d",
X"4a",
X"03",
X"20",
X"56",
X"e4",
X"10",
X"03",
X"4c",
X"25",
X"f1",
X"e8",
X"d0",
X"fd",
X"c8",
X"10",
X"fa",
X"20",
X"b2",
X"f3",
X"a5",
X"06",
X"05",
X"07",
X"f0",
X"12",
X"a5",
X"06",
X"f0",
X"03",
X"ad",
X"fd",
X"bf",
X"a6",
X"07",
X"f0",
X"03",
X"0d",
X"fd",
X"9f",
X"29",
X"01",
X"f0",
X"03",
X"20",
X"cf",
X"f2",
X"a9",
X"00",
X"8d",
X"44",
X"02",
X"a5",
X"06",
X"f0",
X"0a",
X"ad",
X"fd",
X"bf",
X"29",
X"04",
X"f0",
X"03",
X"6c",
X"fa",
X"bf",
X"a5",
X"07",
X"f0",
X"0a",
X"ad",
X"fd",
X"9f",
X"29",
X"04",
X"f0",
X"df",
X"6c",
X"fa",
X"9f",
X"6c",
X"0a",
X"00",
X"a2",
X"f2",
X"a0",
X"f0",
X"20",
X"85",
X"f3",
X"20",
X"30",
X"f2",
X"4c",
X"2a",
X"f2",
X"ad",
X"05",
X"e4",
X"48",
X"ad",
X"04",
X"e4",
X"48",
X"60",
X"6c",
X"fe",
X"bf",
X"6c",
X"fe",
X"9f",
X"c9",
X"d0",
X"d0",
X"1c",
X"60",
X"ee",
X"fc",
X"bf",
X"ad",
X"fc",
X"bf",
X"d0",
X"08",
X"ad",
X"fd",
X"bf",
X"10",
X"03",
X"6c",
X"fe",
X"bf",
X"ce",
X"fc",
X"bf",
X"a0",
X"00",
X"84",
X"05",
X"a9",
X"10",
X"85",
X"06",
X"b1",
X"05",
X"49",
X"ff",
X"91",
X"05",
X"d1",
X"05",
X"d0",
X"da",
X"49",
X"ff",
X"91",
X"05",
X"a5",
X"06",
X"18",
X"69",
X"10",
X"85",
X"06",
X"4c",
X"3f",
X"f2",
X"a9",
X"00",
X"aa",
X"9d",
X"00",
X"d0",
X"9d",
X"00",
X"d4",
X"9d",
X"00",
X"d2",
X"ea",
X"ea",
X"ea",
X"e8",
X"d0",
X"f1",
X"60",
X"c6",
X"11",
X"a9",
X"54",
X"8d",
X"36",
X"02",
X"a9",
X"e7",
X"8d",
X"37",
X"02",
X"a5",
X"06",
X"8d",
X"e4",
X"02",
X"8d",
X"e6",
X"02",
X"a9",
X"00",
X"8d",
X"e5",
X"02",
X"a9",
X"00",
X"8d",
X"e7",
X"02",
X"a9",
X"07",
X"8d",
X"e8",
X"02",
X"20",
X"0c",
X"e4",
X"20",
X"1c",
X"e4",
X"20",
X"2c",
X"e4",
X"20",
X"3c",
X"e4",
X"20",
X"4c",
X"e4",
X"20",
X"6e",
X"e4",
X"20",
X"65",
X"e4",
X"20",
X"6b",
X"e4",
X"ad",
X"1f",
X"d0",
X"29",
X"01",
X"d0",
X"02",
X"e6",
X"4a",
X"60",
X"a5",
X"08",
X"f0",
X"0a",
X"a5",
X"09",
X"29",
X"01",
X"f0",
X"03",
X"20",
X"7e",
X"f3",
X"60",
X"a9",
X"01",
X"8d",
X"01",
X"03",
X"a9",
X"53",
X"8d",
X"02",
X"03",
X"20",
X"53",
X"e4",
X"10",
X"01",
X"60",
X"a9",
X"00",
X"8d",
X"0b",
X"03",
X"a9",
X"01",
X"8d",
X"0a",
X"03",
X"a9",
X"00",
X"8d",
X"04",
X"03",
X"a9",
X"04",
X"8d",
X"05",
X"03",
X"20",
X"9d",
X"f3",
X"10",
X"08",
X"20",
X"81",
X"f3",
X"a5",
X"4b",
X"f0",
X"e0",
X"60",
X"a2",
X"03",
X"bd",
X"00",
X"04",
X"9d",
X"40",
X"02",
X"ca",
X"10",
X"f7",
X"ad",
X"42",
X"02",
X"85",
X"04",
X"ad",
X"43",
X"02",
X"85",
X"05",
X"ad",
X"04",
X"04",
X"85",
X"0c",
X"ad",
X"05",
X"04",
X"85",
X"0d",
X"a0",
X"7f",
X"b9",
X"00",
X"04",
X"91",
X"04",
X"88",
X"10",
X"f8",
X"18",
X"a5",
X"04",
X"69",
X"80",
X"85",
X"04",
X"a5",
X"05",
X"69",
X"00",
X"85",
X"05",
X"ce",
X"41",
X"02",
X"f0",
X"11",
X"ee",
X"0a",
X"03",
X"20",
X"9d",
X"f3",
X"10",
X"dc",
X"20",
X"81",
X"f3",
X"a5",
X"4b",
X"d0",
X"ae",
X"f0",
X"f2",
X"a5",
X"4b",
X"f0",
X"03",
X"20",
X"9d",
X"f3",
X"20",
X"6c",
X"f3",
X"b0",
X"a0",
X"20",
X"7e",
X"f3",
X"e6",
X"09",
X"60",
X"18",
X"ad",
X"42",
X"02",
X"69",
X"06",
X"85",
X"04",
X"ad",
X"43",
X"02",
X"69",
X"00",
X"85",
X"05",
X"6c",
X"04",
X"00",
X"6c",
X"0c",
X"00",
X"a2",
X"0d",
X"a0",
X"f1",
X"8a",
X"a2",
X"00",
X"9d",
X"44",
X"03",
X"98",
X"9d",
X"45",
X"03",
X"a9",
X"09",
X"9d",
X"42",
X"03",
X"a9",
X"ff",
X"9d",
X"48",
X"03",
X"20",
X"56",
X"e4",
X"60",
X"a5",
X"4b",
X"f0",
X"03",
X"4c",
X"7a",
X"e4",
X"a9",
X"52",
X"8d",
X"02",
X"03",
X"a9",
X"01",
X"8d",
X"01",
X"03",
X"20",
X"53",
X"e4",
X"60",
X"a5",
X"08",
X"f0",
X"0a",
X"a5",
X"09",
X"29",
X"02",
X"f0",
X"03",
X"20",
X"e1",
X"f3",
X"60",
X"a5",
X"4a",
X"f0",
X"1c",
X"a9",
X"80",
X"85",
X"3e",
X"e6",
X"4b",
X"20",
X"7d",
X"e4",
X"20",
X"01",
X"f3",
X"a9",
X"00",
X"85",
X"4b",
X"85",
X"4a",
X"06",
X"09",
X"a5",
X"0c",
X"85",
X"02",
X"a5",
X"0d",
X"85",
X"03",
X"60",
X"6c",
X"02",
X"00",
X"a9",
X"ff",
X"8d",
X"fc",
X"02",
X"ad",
X"e6",
X"02",
X"29",
X"f0",
X"85",
X"6a",
X"a9",
X"40",
X"8d",
X"be",
X"02",
X"60",
X"a5",
X"2b",
X"29",
X"0f",
X"d0",
X"08",
X"a5",
X"2a",
X"29",
X"0f",
X"85",
X"2a",
X"a9",
X"00",
X"85",
X"57",
X"a9",
X"e0",
X"8d",
X"f4",
X"02",
X"a9",
X"02",
X"8d",
X"f3",
X"02",
X"8d",
X"2f",
X"02",
X"a9",
X"01",
X"85",
X"4c",
X"a9",
X"c0",
X"05",
X"10",
X"85",
X"10",
X"8d",
X"0e",
X"d2",
X"a9",
X"00",
X"8d",
X"93",
X"02",
X"85",
X"64",
X"85",
X"7b",
X"8d",
X"f0",
X"02",
X"a0",
X"0e",
X"a9",
X"01",
X"99",
X"a3",
X"02",
X"88",
X"10",
X"fa",
X"a2",
X"04",
X"bd",
X"c1",
X"fe",
X"9d",
X"c4",
X"02",
X"ca",
X"10",
X"f7",
X"a4",
X"6a",
X"88",
X"8c",
X"95",
X"02",
X"a9",
X"60",
X"8d",
X"94",
X"02",
X"a6",
X"57",
X"bd",
X"69",
X"fe",
X"d0",
X"04",
X"a9",
X"91",
X"85",
X"4c",
X"85",
X"51",
X"a5",
X"6a",
X"85",
X"65",
X"bc",
X"45",
X"fe",
X"a9",
X"28",
X"20",
X"21",
X"f9",
X"88",
X"d0",
X"f8",
X"ad",
X"6f",
X"02",
X"29",
X"3f",
X"85",
X"67",
X"a8",
X"e0",
X"08",
X"90",
X"17",
X"8a",
X"6a",
X"6a",
X"6a",
X"29",
X"c0",
X"05",
X"67",
X"a8",
X"a9",
X"10",
X"20",
X"21",
X"f9",
X"e0",
X"0b",
X"d0",
X"05",
X"a9",
X"06",
X"8d",
X"c8",
X"02",
X"8c",
X"6f",
X"02",
X"a5",
X"64",
X"85",
X"58",
X"a5",
X"65",
X"85",
X"59",
X"ad",
X"0b",
X"d4",
X"c9",
X"7a",
X"d0",
X"f9",
X"20",
X"1f",
X"f9",
X"bd",
X"75",
X"fe",
X"f0",
X"06",
X"a9",
X"ff",
X"85",
X"64",
X"c6",
X"65",
X"a5",
X"64",
X"85",
X"68",
X"a5",
X"65",
X"85",
X"69",
X"20",
X"13",
X"f9",
X"a9",
X"41",
X"20",
X"17",
X"f9",
X"86",
X"66",
X"a9",
X"18",
X"8d",
X"bf",
X"02",
X"a5",
X"57",
X"c9",
X"09",
X"b0",
X"2d",
X"a5",
X"2a",
X"29",
X"10",
X"f0",
X"27",
X"a9",
X"04",
X"8d",
X"bf",
X"02",
X"a2",
X"02",
X"a9",
X"02",
X"20",
X"17",
X"f9",
X"ca",
X"10",
X"f8",
X"a4",
X"6a",
X"88",
X"98",
X"20",
X"17",
X"f9",
X"a9",
X"60",
X"20",
X"17",
X"f9",
X"a9",
X"42",
X"20",
X"17",
X"f9",
X"18",
X"a9",
X"0c",
X"65",
X"66",
X"85",
X"66",
X"a4",
X"66",
X"be",
X"51",
X"fe",
X"a5",
X"51",
X"20",
X"17",
X"f9",
X"ca",
X"d0",
X"f8",
X"a5",
X"57",
X"c9",
X"08",
X"90",
X"1c",
X"a2",
X"5d",
X"a5",
X"6a",
X"38",
X"e9",
X"10",
X"20",
X"17",
X"f9",
X"a9",
X"00",
X"20",
X"17",
X"f9",
X"a9",
X"4f",
X"20",
X"17",
X"f9",
X"a5",
X"51",
X"20",
X"17",
X"f9",
X"ca",
X"d0",
X"f8",
X"a5",
X"59",
X"20",
X"17",
X"f9",
X"a5",
X"58",
X"20",
X"17",
X"f9",
X"a5",
X"51",
X"09",
X"40",
X"20",
X"17",
X"f9",
X"a9",
X"70",
X"20",
X"17",
X"f9",
X"a9",
X"70",
X"20",
X"17",
X"f9",
X"a5",
X"64",
X"8d",
X"30",
X"02",
X"a5",
X"65",
X"8d",
X"31",
X"02",
X"a9",
X"70",
X"20",
X"17",
X"f9",
X"a5",
X"64",
X"8d",
X"e5",
X"02",
X"a5",
X"65",
X"8d",
X"e6",
X"02",
X"a5",
X"68",
X"85",
X"64",
X"a5",
X"69",
X"85",
X"65",
X"ad",
X"31",
X"02",
X"20",
X"17",
X"f9",
X"ad",
X"30",
X"02",
X"20",
X"17",
X"f9",
X"a5",
X"4c",
X"10",
X"07",
X"48",
X"20",
X"fc",
X"f3",
X"68",
X"a8",
X"60",
X"a5",
X"2a",
X"29",
X"20",
X"d0",
X"0b",
X"20",
X"b9",
X"f7",
X"8d",
X"90",
X"02",
X"a5",
X"52",
X"8d",
X"91",
X"02",
X"a9",
X"22",
X"0d",
X"2f",
X"02",
X"8d",
X"2f",
X"02",
X"4c",
X"21",
X"f6",
X"20",
X"96",
X"fa",
X"20",
X"a2",
X"f5",
X"20",
X"32",
X"fb",
X"20",
X"d4",
X"f9",
X"4c",
X"34",
X"f6",
X"20",
X"47",
X"f9",
X"b1",
X"64",
X"2d",
X"a0",
X"02",
X"46",
X"6f",
X"b0",
X"03",
X"4a",
X"10",
X"f9",
X"8d",
X"fa",
X"02",
X"c9",
X"00",
X"60",
X"8d",
X"fb",
X"02",
X"20",
X"96",
X"fa",
X"ad",
X"fb",
X"02",
X"c9",
X"7d",
X"d0",
X"06",
X"20",
X"b9",
X"f7",
X"4c",
X"21",
X"f6",
X"ad",
X"fb",
X"02",
X"c9",
X"9b",
X"d0",
X"06",
X"20",
X"30",
X"fa",
X"4c",
X"21",
X"f6",
X"20",
X"e0",
X"f5",
X"20",
X"d8",
X"f9",
X"4c",
X"21",
X"f6",
X"ad",
X"ff",
X"02",
X"d0",
X"fb",
X"a2",
X"02",
X"b5",
X"54",
X"95",
X"5a",
X"ca",
X"10",
X"f9",
X"ad",
X"fb",
X"02",
X"a8",
X"2a",
X"2a",
X"2a",
X"2a",
X"29",
X"03",
X"aa",
X"98",
X"29",
X"9f",
X"1d",
X"f6",
X"fe",
X"8d",
X"fa",
X"02",
X"20",
X"47",
X"f9",
X"ad",
X"fa",
X"02",
X"46",
X"6f",
X"b0",
X"04",
X"0a",
X"4c",
X"08",
X"f6",
X"2d",
X"a0",
X"02",
X"85",
X"50",
X"ad",
X"a0",
X"02",
X"49",
X"ff",
X"31",
X"64",
X"05",
X"50",
X"91",
X"64",
X"60",
X"20",
X"a2",
X"f5",
X"85",
X"5d",
X"a6",
X"57",
X"d0",
X"0a",
X"ae",
X"f0",
X"02",
X"d0",
X"05",
X"49",
X"80",
X"20",
X"ff",
X"f5",
X"a4",
X"4c",
X"a9",
X"01",
X"85",
X"4c",
X"ad",
X"fb",
X"02",
X"60",
X"20",
X"b3",
X"fc",
X"20",
X"88",
X"fa",
X"a5",
X"6b",
X"d0",
X"34",
X"a5",
X"54",
X"85",
X"6c",
X"a5",
X"55",
X"85",
X"6d",
X"20",
X"e2",
X"f6",
X"84",
X"4c",
X"ad",
X"fb",
X"02",
X"c9",
X"9b",
X"f0",
X"12",
X"20",
X"ad",
X"f6",
X"20",
X"b3",
X"fc",
X"a5",
X"63",
X"c9",
X"71",
X"d0",
X"03",
X"20",
X"0a",
X"f9",
X"4c",
X"50",
X"f6",
X"20",
X"e4",
X"fa",
X"20",
X"00",
X"fc",
X"a5",
X"6c",
X"85",
X"54",
X"a5",
X"6d",
X"85",
X"55",
X"a5",
X"6b",
X"f0",
X"11",
X"c6",
X"6b",
X"f0",
X"0d",
X"a5",
X"4c",
X"30",
X"f8",
X"20",
X"93",
X"f5",
X"8d",
X"fb",
X"02",
X"4c",
X"b3",
X"fc",
X"20",
X"30",
X"fa",
X"a9",
X"9b",
X"8d",
X"fb",
X"02",
X"20",
X"21",
X"f6",
X"84",
X"4c",
X"4c",
X"b3",
X"fc",
X"6c",
X"64",
X"00",
X"8d",
X"fb",
X"02",
X"20",
X"b3",
X"fc",
X"20",
X"88",
X"fa",
X"20",
X"e4",
X"fa",
X"20",
X"8d",
X"fc",
X"f0",
X"09",
X"0e",
X"a2",
X"02",
X"20",
X"ca",
X"f5",
X"4c",
X"b3",
X"fc",
X"ad",
X"fe",
X"02",
X"0d",
X"a2",
X"02",
X"d0",
X"ef",
X"0e",
X"a2",
X"02",
X"e8",
X"bd",
X"c6",
X"fe",
X"85",
X"64",
X"bd",
X"c7",
X"fe",
X"85",
X"65",
X"20",
X"a1",
X"f6",
X"20",
X"21",
X"f6",
X"4c",
X"b3",
X"fc",
X"a9",
X"ff",
X"8d",
X"fc",
X"02",
X"a5",
X"2a",
X"4a",
X"b0",
X"62",
X"a9",
X"80",
X"a6",
X"11",
X"f0",
X"58",
X"ad",
X"fc",
X"02",
X"c9",
X"ff",
X"f0",
X"ee",
X"85",
X"7c",
X"a2",
X"ff",
X"8e",
X"fc",
X"02",
X"20",
X"d8",
X"fc",
X"aa",
X"e0",
X"c0",
X"90",
X"02",
X"a2",
X"03",
X"bd",
X"fe",
X"fe",
X"8d",
X"fb",
X"02",
X"c9",
X"80",
X"f0",
X"ce",
X"c9",
X"81",
X"d0",
X"0b",
X"ad",
X"b6",
X"02",
X"49",
X"80",
X"8d",
X"b6",
X"02",
X"4c",
X"dd",
X"f6",
X"c9",
X"82",
X"d0",
X"07",
X"a9",
X"00",
X"8d",
X"be",
X"02",
X"f0",
X"b4",
X"c9",
X"83",
X"d0",
X"07",
X"a9",
X"40",
X"8d",
X"be",
X"02",
X"d0",
X"a9",
X"c9",
X"84",
X"d0",
X"07",
X"a9",
X"80",
X"8d",
X"be",
X"02",
X"d0",
X"9e",
X"c9",
X"85",
X"d0",
X"0a",
X"a9",
X"88",
X"85",
X"4c",
X"85",
X"11",
X"a9",
X"9b",
X"d0",
X"26",
X"a5",
X"7c",
X"c9",
X"40",
X"b0",
X"15",
X"ad",
X"fb",
X"02",
X"c9",
X"61",
X"90",
X"0e",
X"c9",
X"7b",
X"b0",
X"0a",
X"ad",
X"be",
X"02",
X"f0",
X"05",
X"05",
X"7c",
X"4c",
X"fe",
X"f6",
X"20",
X"8d",
X"fc",
X"f0",
X"09",
X"ad",
X"fb",
X"02",
X"4d",
X"b6",
X"02",
X"8d",
X"fb",
X"02",
X"4c",
X"34",
X"f6",
X"a9",
X"80",
X"8d",
X"a2",
X"02",
X"60",
X"c6",
X"54",
X"10",
X"06",
X"ae",
X"bf",
X"02",
X"ca",
X"86",
X"54",
X"4c",
X"5c",
X"fc",
X"e6",
X"54",
X"a5",
X"54",
X"cd",
X"bf",
X"02",
X"90",
X"f4",
X"a2",
X"00",
X"f0",
X"ee",
X"c6",
X"55",
X"a5",
X"55",
X"30",
X"04",
X"c5",
X"52",
X"b0",
X"04",
X"a5",
X"53",
X"85",
X"55",
X"4c",
X"dd",
X"fb",
X"e6",
X"55",
X"a5",
X"55",
X"c5",
X"53",
X"90",
X"f5",
X"f0",
X"f3",
X"a5",
X"52",
X"4c",
X"a5",
X"f7",
X"20",
X"f3",
X"fc",
X"a0",
X"00",
X"98",
X"91",
X"64",
X"c8",
X"d0",
X"fb",
X"e6",
X"65",
X"a6",
X"65",
X"e4",
X"6a",
X"90",
X"f3",
X"a9",
X"ff",
X"99",
X"b2",
X"02",
X"c8",
X"c0",
X"04",
X"90",
X"f8",
X"20",
X"e4",
X"fc",
X"85",
X"63",
X"85",
X"6d",
X"a9",
X"00",
X"85",
X"54",
X"85",
X"56",
X"85",
X"6c",
X"60",
X"a5",
X"63",
X"c5",
X"52",
X"f0",
X"21",
X"a5",
X"55",
X"c5",
X"52",
X"d0",
X"03",
X"20",
X"73",
X"fc",
X"20",
X"99",
X"f7",
X"a5",
X"55",
X"c5",
X"53",
X"d0",
X"07",
X"a5",
X"54",
X"f0",
X"03",
X"20",
X"7f",
X"f7",
X"a9",
X"20",
X"8d",
X"fb",
X"02",
X"20",
X"e0",
X"f5",
X"4c",
X"dd",
X"fb",
X"20",
X"aa",
X"f7",
X"a5",
X"55",
X"c5",
X"52",
X"d0",
X"0a",
X"20",
X"34",
X"fa",
X"20",
X"20",
X"fb",
X"90",
X"02",
X"b0",
X"07",
X"a5",
X"63",
X"20",
X"25",
X"fb",
X"90",
X"e6",
X"4c",
X"dd",
X"fb",
X"a5",
X"63",
X"4c",
X"06",
X"fb",
X"a5",
X"63",
X"4c",
X"12",
X"fb",
X"20",
X"9d",
X"fc",
X"20",
X"a2",
X"f5",
X"85",
X"7d",
X"a9",
X"00",
X"8d",
X"bb",
X"02",
X"20",
X"ff",
X"f5",
X"a5",
X"63",
X"48",
X"20",
X"dc",
X"f9",
X"68",
X"c5",
X"63",
X"b0",
X"0c",
X"a5",
X"7d",
X"48",
X"20",
X"a2",
X"f5",
X"85",
X"7d",
X"68",
X"4c",
X"44",
X"f8",
X"20",
X"a8",
X"fc",
X"ce",
X"bb",
X"02",
X"30",
X"04",
X"c6",
X"54",
X"d0",
X"f7",
X"4c",
X"dd",
X"fb",
X"20",
X"9d",
X"fc",
X"20",
X"47",
X"f9",
X"a5",
X"64",
X"85",
X"68",
X"a5",
X"65",
X"85",
X"69",
X"a5",
X"63",
X"48",
X"20",
X"d4",
X"f9",
X"68",
X"c5",
X"63",
X"b0",
X"10",
X"a5",
X"54",
X"cd",
X"bf",
X"02",
X"b0",
X"09",
X"20",
X"a2",
X"f5",
X"a0",
X"00",
X"91",
X"68",
X"f0",
X"da",
X"a0",
X"00",
X"98",
X"91",
X"68",
X"20",
X"68",
X"fc",
X"20",
X"a8",
X"fc",
X"4c",
X"dd",
X"fb",
X"38",
X"20",
X"7b",
X"fb",
X"a5",
X"52",
X"85",
X"55",
X"20",
X"47",
X"f9",
X"a5",
X"64",
X"85",
X"68",
X"18",
X"69",
X"28",
X"85",
X"66",
X"a5",
X"65",
X"85",
X"69",
X"69",
X"00",
X"85",
X"67",
X"a6",
X"54",
X"e0",
X"17",
X"f0",
X"08",
X"20",
X"4e",
X"fb",
X"e8",
X"e0",
X"17",
X"d0",
X"f8",
X"20",
X"9b",
X"fb",
X"4c",
X"dd",
X"fb",
X"20",
X"dd",
X"fb",
X"a4",
X"51",
X"84",
X"54",
X"a4",
X"54",
X"98",
X"38",
X"20",
X"23",
X"fb",
X"08",
X"98",
X"18",
X"69",
X"78",
X"28",
X"20",
X"04",
X"fb",
X"c8",
X"c0",
X"18",
X"d0",
X"ed",
X"ad",
X"b4",
X"02",
X"09",
X"01",
X"8d",
X"b4",
X"02",
X"a5",
X"52",
X"85",
X"55",
X"20",
X"47",
X"f9",
X"20",
X"b7",
X"fb",
X"20",
X"20",
X"fb",
X"90",
X"d4",
X"4c",
X"dd",
X"fb",
X"60",
X"20",
X"20",
X"d8",
X"fc",
X"88",
X"10",
X"fa",
X"60",
X"a9",
X"02",
X"d0",
X"0a",
X"a4",
X"4c",
X"30",
X"2b",
X"a0",
X"00",
X"91",
X"64",
X"a9",
X"01",
X"8d",
X"9e",
X"02",
X"a5",
X"4c",
X"30",
X"1e",
X"a5",
X"64",
X"38",
X"ed",
X"9e",
X"02",
X"85",
X"64",
X"b0",
X"02",
X"c6",
X"65",
X"a5",
X"0f",
X"c5",
X"65",
X"90",
X"0c",
X"d0",
X"06",
X"a5",
X"0e",
X"c5",
X"64",
X"90",
X"04",
X"a9",
X"93",
X"85",
X"4c",
X"60",
X"a5",
X"54",
X"48",
X"a5",
X"55",
X"48",
X"a5",
X"56",
X"48",
X"20",
X"f3",
X"fc",
X"a5",
X"54",
X"85",
X"66",
X"a9",
X"00",
X"85",
X"67",
X"a5",
X"66",
X"0a",
X"26",
X"67",
X"85",
X"51",
X"a4",
X"67",
X"8c",
X"9f",
X"02",
X"0a",
X"26",
X"67",
X"0a",
X"26",
X"67",
X"18",
X"65",
X"51",
X"85",
X"66",
X"a5",
X"67",
X"6d",
X"9f",
X"02",
X"85",
X"67",
X"a6",
X"57",
X"bc",
X"81",
X"fe",
X"88",
X"30",
X"07",
X"06",
X"66",
X"26",
X"67",
X"4c",
X"7e",
X"f9",
X"bc",
X"a5",
X"fe",
X"a5",
X"55",
X"a2",
X"07",
X"88",
X"30",
X"0a",
X"ca",
X"46",
X"56",
X"6a",
X"6e",
X"a1",
X"02",
X"4c",
X"8f",
X"f9",
X"c8",
X"18",
X"65",
X"66",
X"85",
X"66",
X"90",
X"02",
X"e6",
X"67",
X"38",
X"6e",
X"a1",
X"02",
X"18",
X"ca",
X"10",
X"f9",
X"ae",
X"a1",
X"02",
X"a5",
X"66",
X"18",
X"65",
X"64",
X"85",
X"64",
X"85",
X"5e",
X"a5",
X"67",
X"65",
X"65",
X"85",
X"65",
X"85",
X"5f",
X"bd",
X"b1",
X"fe",
X"8d",
X"a0",
X"02",
X"85",
X"6f",
X"68",
X"85",
X"56",
X"68",
X"85",
X"55",
X"68",
X"85",
X"54",
X"60",
X"a9",
X"00",
X"f0",
X"02",
X"a9",
X"9b",
X"85",
X"7d",
X"e6",
X"63",
X"e6",
X"55",
X"d0",
X"02",
X"e6",
X"56",
X"a5",
X"55",
X"a6",
X"57",
X"dd",
X"8d",
X"fe",
X"f0",
X"0b",
X"e0",
X"00",
X"d0",
X"06",
X"c5",
X"53",
X"f0",
X"02",
X"b0",
X"01",
X"60",
X"e0",
X"08",
X"90",
X"04",
X"a5",
X"56",
X"f0",
X"f7",
X"a5",
X"57",
X"d0",
X"30",
X"a5",
X"63",
X"c9",
X"51",
X"90",
X"0a",
X"a5",
X"7d",
X"f0",
X"26",
X"20",
X"30",
X"fa",
X"4c",
X"77",
X"fa",
X"20",
X"34",
X"fa",
X"a5",
X"54",
X"18",
X"69",
X"78",
X"20",
X"25",
X"fb",
X"90",
X"08",
X"a5",
X"7d",
X"f0",
X"04",
X"18",
X"20",
X"a5",
X"f8",
X"4c",
X"dd",
X"fb",
X"a9",
X"00",
X"f0",
X"02",
X"a9",
X"9b",
X"85",
X"7d",
X"20",
X"e4",
X"fc",
X"a9",
X"00",
X"85",
X"56",
X"e6",
X"54",
X"a6",
X"57",
X"a0",
X"18",
X"24",
X"7b",
X"10",
X"05",
X"a0",
X"04",
X"98",
X"d0",
X"03",
X"bd",
X"99",
X"fe",
X"c5",
X"54",
X"d0",
X"26",
X"8c",
X"9d",
X"02",
X"8a",
X"d0",
X"20",
X"a5",
X"7d",
X"f0",
X"1c",
X"c9",
X"9b",
X"38",
X"f0",
X"01",
X"18",
X"20",
X"ac",
X"fb",
X"ee",
X"bb",
X"02",
X"c6",
X"6c",
X"ce",
X"9d",
X"02",
X"ad",
X"b2",
X"02",
X"38",
X"10",
X"ef",
X"ad",
X"9d",
X"02",
X"85",
X"54",
X"4c",
X"dd",
X"fb",
X"38",
X"b5",
X"70",
X"e5",
X"74",
X"95",
X"70",
X"b5",
X"71",
X"e5",
X"75",
X"95",
X"71",
X"60",
X"ad",
X"bf",
X"02",
X"c9",
X"04",
X"f0",
X"07",
X"a5",
X"57",
X"f0",
X"03",
X"20",
X"fc",
X"f3",
X"a9",
X"27",
X"c5",
X"53",
X"b0",
X"02",
X"85",
X"53",
X"a6",
X"57",
X"bd",
X"99",
X"fe",
X"c5",
X"54",
X"90",
X"2a",
X"f0",
X"28",
X"e0",
X"08",
X"d0",
X"0a",
X"a5",
X"56",
X"f0",
X"13",
X"c9",
X"01",
X"d0",
X"1c",
X"f0",
X"04",
X"a5",
X"56",
X"d0",
X"16",
X"bd",
X"8d",
X"fe",
X"c5",
X"55",
X"90",
X"0f",
X"f0",
X"0d",
X"a9",
X"01",
X"85",
X"4c",
X"a9",
X"80",
X"a6",
X"11",
X"85",
X"11",
X"f0",
X"06",
X"60",
X"20",
X"d6",
X"f7",
X"a9",
X"8d",
X"85",
X"4c",
X"68",
X"68",
X"a5",
X"7b",
X"10",
X"03",
X"20",
X"b9",
X"fc",
X"4c",
X"34",
X"f6",
X"a0",
X"00",
X"a5",
X"5d",
X"91",
X"5e",
X"60",
X"48",
X"29",
X"07",
X"aa",
X"bd",
X"b9",
X"fe",
X"85",
X"6e",
X"68",
X"4a",
X"4a",
X"4a",
X"aa",
X"60",
X"2e",
X"b4",
X"02",
X"2e",
X"b3",
X"02",
X"2e",
X"b2",
X"02",
X"60",
X"90",
X"0c",
X"20",
X"eb",
X"fa",
X"bd",
X"a3",
X"02",
X"05",
X"6e",
X"9d",
X"a3",
X"02",
X"60",
X"20",
X"eb",
X"fa",
X"a5",
X"6e",
X"49",
X"ff",
X"3d",
X"a3",
X"02",
X"9d",
X"a3",
X"02",
X"60",
X"a5",
X"54",
X"18",
X"69",
X"78",
X"20",
X"eb",
X"fa",
X"18",
X"bd",
X"a3",
X"02",
X"25",
X"6e",
X"f0",
X"01",
X"38",
X"60",
X"ad",
X"fa",
X"02",
X"a4",
X"57",
X"c0",
X"03",
X"b0",
X"0f",
X"2a",
X"2a",
X"2a",
X"2a",
X"29",
X"03",
X"aa",
X"ad",
X"fa",
X"02",
X"29",
X"9f",
X"1d",
X"fa",
X"fe",
X"8d",
X"fb",
X"02",
X"60",
X"a9",
X"02",
X"85",
X"65",
X"a9",
X"47",
X"85",
X"64",
X"a0",
X"27",
X"b1",
X"66",
X"85",
X"50",
X"b1",
X"68",
X"91",
X"66",
X"a5",
X"50",
X"91",
X"64",
X"88",
X"10",
X"f1",
X"a5",
X"65",
X"85",
X"69",
X"a5",
X"64",
X"85",
X"68",
X"18",
X"a5",
X"66",
X"69",
X"28",
X"85",
X"66",
X"90",
X"02",
X"e6",
X"67",
X"60",
X"08",
X"a0",
X"17",
X"98",
X"20",
X"22",
X"fb",
X"08",
X"98",
X"18",
X"69",
X"79",
X"28",
X"20",
X"04",
X"fb",
X"88",
X"30",
X"04",
X"c4",
X"54",
X"b0",
X"ec",
X"a5",
X"54",
X"18",
X"69",
X"78",
X"28",
X"4c",
X"04",
X"fb",
X"a5",
X"52",
X"85",
X"55",
X"20",
X"47",
X"f9",
X"a0",
X"27",
X"a9",
X"00",
X"91",
X"64",
X"88",
X"10",
X"fb",
X"60",
X"20",
X"fa",
X"fa",
X"a5",
X"58",
X"85",
X"64",
X"a5",
X"59",
X"85",
X"65",
X"a0",
X"28",
X"b1",
X"64",
X"a6",
X"6a",
X"ca",
X"e4",
X"65",
X"d0",
X"08",
X"a2",
X"d7",
X"e4",
X"64",
X"b0",
X"02",
X"a9",
X"00",
X"a0",
X"00",
X"91",
X"64",
X"e6",
X"64",
X"d0",
X"e5",
X"e6",
X"65",
X"a5",
X"65",
X"c5",
X"6a",
X"d0",
X"dd",
X"4c",
X"dd",
X"fb",
X"a9",
X"00",
X"85",
X"63",
X"a5",
X"54",
X"85",
X"51",
X"a5",
X"51",
X"20",
X"22",
X"fb",
X"b0",
X"0c",
X"a5",
X"63",
X"18",
X"69",
X"28",
X"85",
X"63",
X"c6",
X"51",
X"4c",
X"e5",
X"fb",
X"18",
X"a5",
X"63",
X"65",
X"55",
X"85",
X"63",
X"60",
X"20",
X"9d",
X"fc",
X"a5",
X"63",
X"48",
X"a5",
X"6c",
X"85",
X"54",
X"a5",
X"6d",
X"85",
X"55",
X"a9",
X"01",
X"85",
X"6b",
X"a2",
X"17",
X"a5",
X"7b",
X"10",
X"02",
X"a2",
X"03",
X"e4",
X"54",
X"d0",
X"0b",
X"a5",
X"55",
X"c5",
X"53",
X"d0",
X"05",
X"e6",
X"6b",
X"4c",
X"39",
X"fc",
X"20",
X"d4",
X"f9",
X"e6",
X"6b",
X"a5",
X"63",
X"c5",
X"52",
X"d0",
X"de",
X"c6",
X"54",
X"20",
X"99",
X"f7",
X"20",
X"a2",
X"f5",
X"d0",
X"17",
X"c6",
X"6b",
X"a5",
X"63",
X"c5",
X"52",
X"f0",
X"0f",
X"20",
X"99",
X"f7",
X"a5",
X"55",
X"c5",
X"53",
X"d0",
X"02",
X"c6",
X"54",
X"a5",
X"6b",
X"d0",
X"e4",
X"68",
X"85",
X"63",
X"20",
X"a8",
X"fc",
X"60",
X"20",
X"dd",
X"fb",
X"a5",
X"51",
X"85",
X"6c",
X"a5",
X"52",
X"85",
X"6d",
X"60",
X"a5",
X"63",
X"c5",
X"52",
X"d0",
X"02",
X"c6",
X"54",
X"20",
X"dd",
X"fb",
X"a5",
X"63",
X"c5",
X"52",
X"f0",
X"13",
X"20",
X"47",
X"f9",
X"a5",
X"53",
X"38",
X"e5",
X"52",
X"a8",
X"b1",
X"64",
X"d0",
X"06",
X"88",
X"10",
X"f9",
X"4c",
X"db",
X"f8",
X"60",
X"a2",
X"2d",
X"bd",
X"c6",
X"fe",
X"cd",
X"fb",
X"02",
X"f0",
X"05",
X"ca",
X"ca",
X"ca",
X"10",
X"f3",
X"60",
X"a2",
X"02",
X"b5",
X"54",
X"9d",
X"b8",
X"02",
X"ca",
X"10",
X"f8",
X"60",
X"a2",
X"02",
X"bd",
X"b8",
X"02",
X"95",
X"54",
X"ca",
X"10",
X"f8",
X"60",
X"20",
X"b9",
X"fc",
X"4c",
X"34",
X"f6",
X"ad",
X"bf",
X"02",
X"c9",
X"18",
X"f0",
X"17",
X"a2",
X"0b",
X"b5",
X"54",
X"48",
X"bd",
X"90",
X"02",
X"95",
X"54",
X"68",
X"9d",
X"90",
X"02",
X"ca",
X"10",
X"f1",
X"a5",
X"7b",
X"49",
X"ff",
X"85",
X"7b",
X"60",
X"a2",
X"7f",
X"8e",
X"1f",
X"d0",
X"8e",
X"0a",
X"d4",
X"ca",
X"10",
X"f7",
X"60",
X"a9",
X"00",
X"a6",
X"7b",
X"d0",
X"04",
X"a6",
X"57",
X"d0",
X"02",
X"a5",
X"52",
X"85",
X"55",
X"60",
X"a5",
X"58",
X"85",
X"64",
X"a5",
X"59",
X"85",
X"65",
X"60",
X"a2",
X"00",
X"a5",
X"22",
X"c9",
X"11",
X"f0",
X"08",
X"c9",
X"12",
X"f0",
X"03",
X"a0",
X"84",
X"60",
X"e8",
X"8e",
X"b7",
X"02",
X"a5",
X"54",
X"85",
X"60",
X"a5",
X"55",
X"85",
X"61",
X"a5",
X"56",
X"85",
X"62",
X"a9",
X"01",
X"85",
X"79",
X"85",
X"7a",
X"38",
X"a5",
X"60",
X"e5",
X"5a",
X"85",
X"76",
X"b0",
X"0d",
X"a9",
X"ff",
X"85",
X"79",
X"a5",
X"76",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"85",
X"76",
X"38",
X"a5",
X"61",
X"e5",
X"5b",
X"85",
X"77",
X"a5",
X"62",
X"e5",
X"5c",
X"85",
X"78",
X"b0",
X"16",
X"a9",
X"ff",
X"85",
X"7a",
X"a5",
X"77",
X"49",
X"ff",
X"85",
X"77",
X"a5",
X"78",
X"49",
X"ff",
X"85",
X"78",
X"e6",
X"77",
X"d0",
X"02",
X"e6",
X"78",
X"a2",
X"02",
X"a0",
X"00",
X"84",
X"73",
X"98",
X"95",
X"70",
X"b5",
X"5a",
X"95",
X"54",
X"ca",
X"10",
X"f6",
X"a5",
X"77",
X"e8",
X"a8",
X"a5",
X"78",
X"85",
X"7f",
X"85",
X"75",
X"d0",
X"0b",
X"a5",
X"77",
X"c5",
X"76",
X"b0",
X"05",
X"a5",
X"76",
X"a2",
X"02",
X"a8",
X"98",
X"85",
X"7e",
X"85",
X"74",
X"48",
X"a5",
X"75",
X"4a",
X"68",
X"6a",
X"95",
X"70",
X"a5",
X"7e",
X"05",
X"7f",
X"d0",
X"03",
X"4c",
X"42",
X"fe",
X"18",
X"a5",
X"70",
X"65",
X"76",
X"85",
X"70",
X"90",
X"02",
X"e6",
X"71",
X"a5",
X"71",
X"c5",
X"75",
X"90",
X"14",
X"d0",
X"06",
X"a5",
X"70",
X"c5",
X"74",
X"90",
X"0c",
X"18",
X"a5",
X"54",
X"65",
X"79",
X"85",
X"54",
X"a2",
X"00",
X"20",
X"7a",
X"fa",
X"18",
X"a5",
X"72",
X"65",
X"77",
X"85",
X"72",
X"a5",
X"73",
X"65",
X"78",
X"85",
X"73",
X"c5",
X"75",
X"90",
X"27",
X"d0",
X"06",
X"a5",
X"72",
X"c5",
X"74",
X"90",
X"1f",
X"24",
X"7a",
X"10",
X"10",
X"c6",
X"55",
X"a5",
X"55",
X"c9",
X"ff",
X"d0",
X"0e",
X"a5",
X"56",
X"f0",
X"0a",
X"c6",
X"56",
X"10",
X"06",
X"e6",
X"55",
X"d0",
X"02",
X"e6",
X"56",
X"a2",
X"02",
X"20",
X"7a",
X"fa",
X"20",
X"96",
X"fa",
X"20",
X"e0",
X"f5",
X"ad",
X"b7",
X"02",
X"f0",
X"2f",
X"20",
X"9d",
X"fc",
X"ad",
X"fb",
X"02",
X"8d",
X"bc",
X"02",
X"a5",
X"54",
X"48",
X"20",
X"dc",
X"f9",
X"68",
X"85",
X"54",
X"20",
X"96",
X"fa",
X"20",
X"a2",
X"f5",
X"d0",
X"0c",
X"ad",
X"fd",
X"02",
X"8d",
X"fb",
X"02",
X"20",
X"e0",
X"f5",
X"4c",
X"0a",
X"fe",
X"ad",
X"bc",
X"02",
X"8d",
X"fb",
X"02",
X"20",
X"a8",
X"fc",
X"38",
X"a5",
X"7e",
X"e9",
X"01",
X"85",
X"7e",
X"a5",
X"7f",
X"e9",
X"00",
X"85",
X"7f",
X"30",
X"03",
X"4c",
X"90",
X"fd",
X"4c",
X"34",
X"f6",
X"18",
X"10",
X"0a",
X"0a",
X"10",
X"1c",
X"34",
X"64",
X"c4",
X"c4",
X"c4",
X"c4",
X"17",
X"17",
X"0b",
X"17",
X"2f",
X"2f",
X"5f",
X"5f",
X"61",
X"61",
X"61",
X"61",
X"13",
X"13",
X"09",
X"13",
X"27",
X"27",
X"4f",
X"4f",
X"41",
X"41",
X"41",
X"41",
X"02",
X"06",
X"07",
X"08",
X"09",
X"0a",
X"0b",
X"0d",
X"0f",
X"0f",
X"0f",
X"0f",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"02",
X"01",
X"01",
X"00",
X"00",
X"01",
X"01",
X"02",
X"02",
X"02",
X"02",
X"02",
X"28",
X"14",
X"14",
X"28",
X"50",
X"50",
X"a0",
X"a0",
X"40",
X"50",
X"50",
X"50",
X"18",
X"18",
X"0c",
X"18",
X"30",
X"30",
X"60",
X"60",
X"c0",
X"c0",
X"c0",
X"c0",
X"00",
X"00",
X"00",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"01",
X"01",
X"01",
X"00",
X"ff",
X"f0",
X"0f",
X"c0",
X"30",
X"0c",
X"03",
X"80",
X"40",
X"20",
X"10",
X"08",
X"04",
X"02",
X"01",
X"28",
X"ca",
X"94",
X"46",
X"00",
X"1b",
X"79",
X"f7",
X"1c",
X"7f",
X"f7",
X"1d",
X"8c",
X"f7",
X"1e",
X"99",
X"f7",
X"1f",
X"aa",
X"f7",
X"7d",
X"b9",
X"f7",
X"7e",
X"e6",
X"f7",
X"7f",
X"10",
X"f8",
X"9b",
X"30",
X"fa",
X"9c",
X"d4",
X"f8",
X"9d",
X"a4",
X"f8",
X"9e",
X"32",
X"f8",
X"9f",
X"2d",
X"f8",
X"fd",
X"0a",
X"f9",
X"fe",
X"6d",
X"f8",
X"ff",
X"37",
X"f8",
X"40",
X"00",
X"20",
X"60",
X"20",
X"40",
X"00",
X"60",
X"6c",
X"6a",
X"3b",
X"80",
X"80",
X"6b",
X"2b",
X"2a",
X"6f",
X"80",
X"70",
X"75",
X"9b",
X"69",
X"2d",
X"3d",
X"76",
X"80",
X"63",
X"80",
X"80",
X"62",
X"78",
X"7a",
X"34",
X"80",
X"33",
X"36",
X"1b",
X"35",
X"32",
X"31",
X"2c",
X"20",
X"2e",
X"6e",
X"80",
X"6d",
X"2f",
X"81",
X"72",
X"80",
X"65",
X"79",
X"7f",
X"74",
X"77",
X"71",
X"39",
X"80",
X"30",
X"37",
X"7e",
X"38",
X"3c",
X"3e",
X"66",
X"68",
X"64",
X"80",
X"82",
X"67",
X"73",
X"61",
X"4c",
X"4a",
X"3a",
X"80",
X"80",
X"4b",
X"5c",
X"5e",
X"4f",
X"80",
X"50",
X"55",
X"9b",
X"49",
X"5f",
X"7c",
X"56",
X"80",
X"43",
X"80",
X"80",
X"42",
X"58",
X"5a",
X"24",
X"80",
X"23",
X"26",
X"1b",
X"25",
X"22",
X"21",
X"5b",
X"20",
X"5d",
X"4e",
X"80",
X"4d",
X"3f",
X"81",
X"52",
X"80",
X"45",
X"59",
X"9f",
X"54",
X"57",
X"51",
X"28",
X"80",
X"29",
X"27",
X"9c",
X"40",
X"7d",
X"9d",
X"46",
X"48",
X"44",
X"80",
X"83",
X"47",
X"53",
X"41",
X"0c",
X"0a",
X"7b",
X"80",
X"80",
X"0b",
X"1e",
X"1f",
X"0f",
X"80",
X"10",
X"15",
X"9b",
X"09",
X"1c",
X"1d",
X"16",
X"80",
X"03",
X"80",
X"80",
X"02",
X"18",
X"1a",
X"80",
X"80",
X"85",
X"80",
X"1b",
X"80",
X"fd",
X"80",
X"00",
X"20",
X"60",
X"0e",
X"80",
X"0d",
X"80",
X"81",
X"12",
X"80",
X"05",
X"19",
X"9e",
X"14",
X"17",
X"11",
X"80",
X"80",
X"80",
X"80",
X"fe",
X"80",
X"7d",
X"ff",
X"06",
X"08",
X"04",
X"80",
X"84",
X"07",
X"13",
X"01",
X"ad",
X"09",
X"d2",
X"cd",
X"f2",
X"02",
X"d0",
X"05",
X"ad",
X"f1",
X"02",
X"d0",
X"20",
X"ad",
X"09",
X"d2",
X"c9",
X"9f",
X"d0",
X"0a",
X"ad",
X"ff",
X"02",
X"49",
X"ff",
X"8d",
X"ff",
X"02",
X"b0",
X"0f",
X"8d",
X"fc",
X"02",
X"8d",
X"f2",
X"02",
X"a9",
X"03",
X"8d",
X"f1",
X"02",
X"a9",
X"00",
X"85",
X"4d",
X"a9",
X"30",
X"8d",
X"2b",
X"02",
X"68",
X"40",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"f3",
X"e6",
X"91",
X"e7",
X"25",
X"f1",
X"f3",
X"e6"

);
        signal rdata:std_logic_vector(7 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
