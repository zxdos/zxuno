library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity yuv_table is
	Port (color	: in  std_logic_vector (5 downto 0);
			y		: out std_logic_vector (5 downto 0);
			u		: out std_logic_vector (5 downto 0);
			v		: out std_logic_vector (5 downto 0));
end yuv_table;

architecture Behavioral of yuv_table is
begin

	process (color)
	begin
		case color is
		when "000000" => y <= "000000";
		when "000001" => y <= "000011";
		when "000010" => y <= "000110";
		when "000011" => y <= "001001";
		when "000100" => y <= "000110";
		when "000101" => y <= "001001";
		when "000110" => y <= "001100";
		when "000111" => y <= "001111";
		when "001000" => y <= "001100";
		when "001001" => y <= "001111";
		when "001010" => y <= "010010";
		when "001011" => y <= "010101";
		when "001100" => y <= "010010";
		when "001101" => y <= "010101";
		when "001110" => y <= "011000";
		when "001111" => y <= "011011";
		when "010000" => y <= "000001";
		when "010001" => y <= "000100";
		when "010010" => y <= "000111";
		when "010011" => y <= "001010";
		when "010100" => y <= "000111";
		when "010101" => y <= "001010";
		when "010110" => y <= "001101";
		when "010111" => y <= "010000";
		when "011000" => y <= "001101";
		when "011001" => y <= "010000";
		when "011010" => y <= "010011";
		when "011011" => y <= "010110";
		when "011100" => y <= "010011";
		when "011101" => y <= "010110";
		when "011110" => y <= "011001";
		when "011111" => y <= "011100";
		when "100000" => y <= "000010";
		when "100001" => y <= "000101";
		when "100010" => y <= "001000";
		when "100011" => y <= "001011";
		when "100100" => y <= "001000";
		when "100101" => y <= "001011";
		when "100110" => y <= "001110";
		when "100111" => y <= "010001";
		when "101000" => y <= "001110";
		when "101001" => y <= "010001";
		when "101010" => y <= "010100";
		when "101011" => y <= "010111";
		when "101100" => y <= "010100";
		when "101101" => y <= "010111";
		when "101110" => y <= "011010";
		when "101111" => y <= "011101";
		when "110000" => y <= "000011";
		when "110001" => y <= "000110";
		when "110010" => y <= "001001";
		when "110011" => y <= "001100";
		when "110100" => y <= "001001";
		when "110101" => y <= "001100";
		when "110110" => y <= "001111";
		when "110111" => y <= "010010";
		when "111000" => y <= "001111";
		when "111001" => y <= "010010";
		when "111010" => y <= "010101";
		when "111011" => y <= "011000";
		when "111100" => y <= "010101";
		when "111101" => y <= "011000";
		when "111110" => y <= "011011";
		when "111111" => y <= "011110";
		when others =>
		end case;
	end process;

	process (color)
	begin
		case color is
		when "000000" => u <= "000000";
		when "000001" => u <= "111111";
		when "000010" => u <= "111101";
		when "000011" => u <= "111100";
		when "000100" => u <= "111101";
		when "000101" => u <= "111100";
		when "000110" => u <= "111010";
		when "000111" => u <= "111001";
		when "001000" => u <= "111010";
		when "001001" => u <= "111001";
		when "001010" => u <= "110111";
		when "001011" => u <= "110110";
		when "001100" => u <= "110111";
		when "001101" => u <= "110110";
		when "001110" => u <= "110100";
		when "001111" => u <= "110011";
		when "010000" => u <= "000100";
		when "010001" => u <= "000011";
		when "010010" => u <= "000001";
		when "010011" => u <= "000000";
		when "010100" => u <= "000001";
		when "010101" => u <= "000000";
		when "010110" => u <= "111111";
		when "010111" => u <= "111101";
		when "011000" => u <= "111111";
		when "011001" => u <= "111101";
		when "011010" => u <= "111100";
		when "011011" => u <= "111010";
		when "011100" => u <= "111100";
		when "011101" => u <= "111010";
		when "011110" => u <= "111001";
		when "011111" => u <= "110111";
		when "100000" => u <= "001001";
		when "100001" => u <= "000111";
		when "100010" => u <= "000110";
		when "100011" => u <= "000100";
		when "100100" => u <= "000110";
		when "100101" => u <= "000100";
		when "100110" => u <= "000011";
		when "100111" => u <= "000001";
		when "101000" => u <= "000011";
		when "101001" => u <= "000001";
		when "101010" => u <= "000000";
		when "101011" => u <= "111111";
		when "101100" => u <= "000000";
		when "101101" => u <= "111111";
		when "101110" => u <= "111101";
		when "101111" => u <= "111100";
		when "110000" => u <= "001101";
		when "110001" => u <= "001100";
		when "110010" => u <= "001010";
		when "110011" => u <= "001001";
		when "110100" => u <= "001010";
		when "110101" => u <= "001001";
		when "110110" => u <= "000111";
		when "110111" => u <= "000110";
		when "111000" => u <= "000111";
		when "111001" => u <= "000110";
		when "111010" => u <= "000100";
		when "111011" => u <= "000011";
		when "111100" => u <= "000100";
		when "111101" => u <= "000011";
		when "111110" => u <= "000001";
		when "111111" => u <= "000000";
		when others =>
		end case;
	end process;

	process (color)
	begin
		case color is
		when "000000" => v <= "000000";
		when "000001" => v <= "000110";
		when "000010" => v <= "001100";
		when "000011" => v <= "010010";
		when "000100" => v <= "111011";
		when "000101" => v <= "000001";
		when "000110" => v <= "000111";
		when "000111" => v <= "001101";
		when "001000" => v <= "110110";
		when "001001" => v <= "111100";
		when "001010" => v <= "000010";
		when "001011" => v <= "001000";
		when "001100" => v <= "110001";
		when "001101" => v <= "110111";
		when "001110" => v <= "111101";
		when "001111" => v <= "000011";
		when "010000" => v <= "111111";
		when "010001" => v <= "000101";
		when "010010" => v <= "001011";
		when "010011" => v <= "010001";
		when "010100" => v <= "111010";
		when "010101" => v <= "000000";
		when "010110" => v <= "000110";
		when "010111" => v <= "001100";
		when "011000" => v <= "110101";
		when "011001" => v <= "111011";
		when "011010" => v <= "000001";
		when "011011" => v <= "000111";
		when "011100" => v <= "110000";
		when "011101" => v <= "110110";
		when "011110" => v <= "111100";
		when "011111" => v <= "000010";
		when "100000" => v <= "111110";
		when "100001" => v <= "000100";
		when "100010" => v <= "001010";
		when "100011" => v <= "010000";
		when "100100" => v <= "111001";
		when "100101" => v <= "111111";
		when "100110" => v <= "000101";
		when "100111" => v <= "001011";
		when "101000" => v <= "110100";
		when "101001" => v <= "111010";
		when "101010" => v <= "000000";
		when "101011" => v <= "000110";
		when "101100" => v <= "101111";
		when "101101" => v <= "110101";
		when "101110" => v <= "111011";
		when "101111" => v <= "000001";
		when "110000" => v <= "111101";
		when "110001" => v <= "000011";
		when "110010" => v <= "001001";
		when "110011" => v <= "001111";
		when "110100" => v <= "111000";
		when "110101" => v <= "111110";
		when "110110" => v <= "000100";
		when "110111" => v <= "001010";
		when "111000" => v <= "110011";
		when "111001" => v <= "111001";
		when "111010" => v <= "111111";
		when "111011" => v <= "000101";
		when "111100" => v <= "101110";
		when "111101" => v <= "110100";
		when "111110" => v <= "111010";
		when "111111" => v <= "000000";
		when others =>
		end case;
	end process;


end Behavioral;

