
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
	X"0b0b0b89",
X"ad040b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"0b0b0b0b",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fd0608",
X"72830609",
X"81058205",
X"832b2a83",
X"ffff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fd0608",
X"83ffff73",
X"83060981",
X"05820583",
X"2b2b0906",
X"7383ffff",
X"0b0b0b0b",
X"83a70400",
X"72098105",
X"72057373",
X"09060906",
X"73097306",
X"070a8106",
X"53510400",
X"00000000",
X"00000000",
X"72722473",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71737109",
X"71068106",
X"30720a10",
X"0a720a10",
X"0a31050a",
X"81065151",
X"53510400",
X"00000000",
X"72722673",
X"732e0753",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"bc040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"720a722b",
X"0a535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72729f06",
X"0981050b",
X"0b0b889f",
X"05040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72722aff",
X"739f062a",
X"0974090a",
X"8106ff05",
X"06075351",
X"04000000",
X"00000000",
X"00000000",
X"71715351",
X"020d0406",
X"73830609",
X"81058205",
X"832b0b2b",
X"0772fc06",
X"0c515104",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a810653",
X"51040000",
X"00000000",
X"00000000",
X"00000000",
X"72098105",
X"72050970",
X"81050906",
X"0a098106",
X"53510400",
X"00000000",
X"00000000",
X"00000000",
X"71098105",
X"52040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72720981",
X"05055351",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097206",
X"73730906",
X"07535104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"71fc0608",
X"72830609",
X"81058305",
X"1010102a",
X"81ff0652",
X"04000000",
X"00000000",
X"00000000",
X"71fc0608",
X"0b0b80f6",
X"b4738306",
X"10100508",
X"060b0b0b",
X"88a20400",
X"00000000",
X"00000000",
X"0b0b0b88",
X"ff040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"0b0b0b88",
X"d8040000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"72097081",
X"0509060a",
X"8106ff05",
X"70547106",
X"73097274",
X"05ff0506",
X"07515151",
X"04000000",
X"72097081",
X"0509060a",
X"098106ff",
X"05705471",
X"06730972",
X"7405ff05",
X"06075151",
X"51040000",
X"05ff0504",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"810b80fa",
X"f80c5104",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007181",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000284",
X"05721010",
X"05520400",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00007171",
X"05ff0571",
X"5351020d",
X"04000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101010",
X"10101053",
X"51047381",
X"ff067383",
X"06098105",
X"83051010",
X"102b0772",
X"fc060c51",
X"51043c04",
X"72728072",
X"8106ff05",
X"09720605",
X"71105272",
X"0a100a53",
X"72ed3851",
X"51535104",
X"83e08008",
X"83e08408",
X"83e08808",
X"757580f3",
X"e32d5050",
X"83e08008",
X"5683e088",
X"0c83e084",
X"0c83e080",
X"0c510483",
X"e0800883",
X"e0840883",
X"e0880875",
X"7580f3a2",
X"2d505083",
X"e0800856",
X"83e0880c",
X"83e0840c",
X"83e0800c",
X"51040000",
X"800489aa",
X"0489aa0b",
X"80ddb104",
X"fd3d0d75",
X"705254ae",
X"a43f83e0",
X"80081453",
X"72742e92",
X"38ff1370",
X"33535371",
X"af2e0981",
X"06ee3881",
X"13537283",
X"e0800c85",
X"3d0d04fd",
X"3d0d7577",
X"70535454",
X"c73f83e0",
X"8008732e",
X"a13883e0",
X"80087331",
X"52ff1252",
X"71ff2e8f",
X"38727081",
X"05543374",
X"70810556",
X"34eb39ff",
X"14548074",
X"34853d0d",
X"04803d0d",
X"7251ff90",
X"3f823d0d",
X"047183e0",
X"800c0480",
X"3d0d7251",
X"80713481",
X"0bbc120c",
X"800b80c0",
X"120c823d",
X"0d04800b",
X"83e2c008",
X"248a38b4",
X"f53fff0b",
X"83e2c00c",
X"800b83e0",
X"800c04ff",
X"3d0d7352",
X"83e09c08",
X"722e8d38",
X"d93f7151",
X"96993f71",
X"83e09c0c",
X"833d0d04",
X"f43d0d7e",
X"60625c5a",
X"558154bc",
X"15088191",
X"387451cf",
X"3f795880",
X"7a2580f7",
X"3883e2f0",
X"0870892a",
X"5783ff06",
X"78848072",
X"31565657",
X"73782583",
X"38735575",
X"83e2c008",
X"2e8438ff",
X"893f83e2",
X"c0088025",
X"a6387589",
X"2b5198dc",
X"3f83e2f0",
X"088f3dfc",
X"11555c54",
X"8152f81b",
X"5196c63f",
X"761483e2",
X"f00c7583",
X"e2c00c74",
X"53765278",
X"51b3a63f",
X"83e08008",
X"83e2f008",
X"1683e2f0",
X"0c787631",
X"761b5b59",
X"56778024",
X"ff8b3861",
X"7a710c54",
X"75547580",
X"2e833881",
X"547383e0",
X"800c8e3d",
X"0d04fc3d",
X"0dfe9b3f",
X"7651feaf",
X"3f863dfc",
X"05537852",
X"775195e9",
X"3f797571",
X"0c5483e0",
X"80085483",
X"e0800880",
X"2e833881",
X"547383e0",
X"800c863d",
X"0d04fe3d",
X"0d7583e2",
X"c0085353",
X"80722489",
X"3871732e",
X"8438fdd6",
X"3f7451fd",
X"ea3f7251",
X"97ae3f83",
X"e0800852",
X"83e08008",
X"802e8338",
X"81527183",
X"e0800c84",
X"3d0d0480",
X"3d0d7280",
X"c0110883",
X"e0800c51",
X"823d0d04",
X"803d0d72",
X"bc110883",
X"e0800c51",
X"823d0d04",
X"80c40b83",
X"e0800c04",
X"fd3d0d75",
X"77715470",
X"535553a9",
X"fc3f82c8",
X"1308bc15",
X"0c82c013",
X"0880c015",
X"0cfceb3f",
X"735193ab",
X"3f7383e0",
X"9c0c83e0",
X"80085383",
X"e0800880",
X"2e833881",
X"537283e0",
X"800c853d",
X"0d04fd3d",
X"0d757755",
X"53fcbf3f",
X"72802ea5",
X"38bc1308",
X"527351a9",
X"863f83e0",
X"80088f38",
X"77527251",
X"ff9a3f83",
X"e0800853",
X"8a3982cc",
X"130853d8",
X"39815372",
X"83e0800c",
X"853d0d04",
X"fe3d0dff",
X"0b83e2c0",
X"0c7483e0",
X"a00c7583",
X"e2bc0caf",
X"da3f83e0",
X"800881ff",
X"06528153",
X"71993883",
X"e2d8518e",
X"943f83e0",
X"80085283",
X"e0800880",
X"2e833872",
X"52715372",
X"83e0800c",
X"843d0d04",
X"fa3d0d78",
X"7a82c412",
X"0882c412",
X"08707224",
X"59565657",
X"5773732e",
X"09810691",
X"3880c016",
X"5280c017",
X"51a6f73f",
X"83e08008",
X"557483e0",
X"800c883d",
X"0d04f63d",
X"0d7c5b80",
X"7b715c54",
X"577a772e",
X"8c38811a",
X"82cc1408",
X"545a72f6",
X"38805980",
X"d9397a54",
X"81578070",
X"7b7b315a",
X"5755ff18",
X"53747325",
X"80c13882",
X"cc140852",
X"7351ff8c",
X"3f800b83",
X"e0800825",
X"a13882cc",
X"140882cc",
X"110882cc",
X"160c7482",
X"cc120c53",
X"75802e86",
X"387282cc",
X"170c7254",
X"80577382",
X"cc150881",
X"17575556",
X"ffb83981",
X"1959800b",
X"ff1b5454",
X"78732583",
X"38815476",
X"81327075",
X"06515372",
X"ff90388c",
X"3d0d04f7",
X"3d0d7b7d",
X"5a5a82d0",
X"5283e2bc",
X"085180e2",
X"a53f83e0",
X"800857f9",
X"e13f7952",
X"83e2c451",
X"95b73f83",
X"e0800854",
X"805383e0",
X"8008732e",
X"09810682",
X"833883e0",
X"a0080b0b",
X"80f7f453",
X"705256a6",
X"b43f0b0b",
X"80f7f452",
X"80c01651",
X"a6a73f75",
X"bc170c73",
X"82c0170c",
X"810b82c4",
X"170c810b",
X"82c8170c",
X"7382cc17",
X"0cff1782",
X"d0175557",
X"81913983",
X"e0ac3370",
X"822a7081",
X"06515455",
X"72818038",
X"74812a81",
X"06587780",
X"f6387484",
X"2a810682",
X"c4150c83",
X"e0ac3381",
X"0682c815",
X"0c795273",
X"51a5ce3f",
X"7351a5e5",
X"3f83e080",
X"081453af",
X"73708105",
X"553472bc",
X"150c83e0",
X"ad527251",
X"a5af3f83",
X"e0a40882",
X"c0150c83",
X"e0ba5280",
X"c01451a5",
X"9c3f7880",
X"2e8d3873",
X"51782d83",
X"e0800880",
X"2e993877",
X"82cc150c",
X"75802e86",
X"387382cc",
X"170c7382",
X"d015ff19",
X"59555676",
X"802e9b38",
X"83e0a452",
X"83e2c451",
X"94ad3f83",
X"e080088a",
X"3883e0ad",
X"335372fe",
X"d2387880",
X"2e893883",
X"e0a00851",
X"fcb83f83",
X"e0a00853",
X"7283e080",
X"0c8b3d0d",
X"04ff3d0d",
X"80527351",
X"fdb53f83",
X"3d0d04f0",
X"3d0d6270",
X"5254f690",
X"3f83e080",
X"08745387",
X"3d705355",
X"55f6b03f",
X"f7903f73",
X"51d33f63",
X"53745283",
X"e0800851",
X"fab83f92",
X"3d0d0471",
X"83e0800c",
X"0480c012",
X"83e0800c",
X"04803d0d",
X"7282c011",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d7282cc",
X"110883e0",
X"800c5182",
X"3d0d0480",
X"3d0d7282",
X"c4110883",
X"e0800c51",
X"823d0d04",
X"f93d0d79",
X"83e09008",
X"57578177",
X"27819638",
X"76881708",
X"27818e38",
X"75335574",
X"822e8938",
X"74832eb3",
X"3880fe39",
X"74547610",
X"83fe0653",
X"76882a8c",
X"17080552",
X"893dfc05",
X"51aa883f",
X"83e08008",
X"80df3802",
X"9d053389",
X"3d337188",
X"2b075656",
X"80d13984",
X"5476822b",
X"83fc0653",
X"76872a8c",
X"17080552",
X"893dfc05",
X"51a9d83f",
X"83e08008",
X"b038029f",
X"05330284",
X"059e0533",
X"71982b71",
X"902b0702",
X"8c059d05",
X"3370882b",
X"72078d3d",
X"337180ff",
X"fffe8006",
X"07515253",
X"57585683",
X"39815574",
X"83e0800c",
X"893d0d04",
X"fb3d0d83",
X"e09008fe",
X"19881208",
X"fe055556",
X"54805674",
X"73278d38",
X"82143375",
X"71299416",
X"08055753",
X"7583e080",
X"0c873d0d",
X"04fc3d0d",
X"7652800b",
X"83e09008",
X"70335152",
X"5370832e",
X"09810691",
X"38951233",
X"94133371",
X"982b7190",
X"2b075555",
X"519b1233",
X"9a133371",
X"882b0774",
X"0783e080",
X"0c55863d",
X"0d04fc3d",
X"0d7683e0",
X"90085555",
X"80752388",
X"15085372",
X"812e8838",
X"88140873",
X"26853881",
X"52b23972",
X"90387333",
X"5271832e",
X"09810685",
X"38901408",
X"53728c16",
X"0c72802e",
X"8d387251",
X"fed63f83",
X"e0800852",
X"85399014",
X"08527190",
X"160c8052",
X"7183e080",
X"0c863d0d",
X"04fa3d0d",
X"7883e090",
X"08712281",
X"057083ff",
X"ff065754",
X"57557380",
X"2e883890",
X"15085372",
X"86388352",
X"80e73973",
X"8f065271",
X"80da3881",
X"1390160c",
X"8c150853",
X"72903883",
X"0b841722",
X"57527376",
X"2780c638",
X"bf398216",
X"33ff0574",
X"842a0652",
X"71b23872",
X"51fcb13f",
X"81527183",
X"e0800827",
X"a8388352",
X"83e08008",
X"88170827",
X"9c3883e0",
X"80088c16",
X"0c83e080",
X"0851fdbc",
X"3f83e080",
X"0890160c",
X"73752380",
X"527183e0",
X"800c883d",
X"0d04f23d",
X"0d606264",
X"585e5b75",
X"335574a0",
X"2e098106",
X"88388116",
X"704456ef",
X"39627033",
X"565674af",
X"2e098106",
X"84388116",
X"43800b88",
X"1c0c6270",
X"33515574",
X"9f269138",
X"7a51fdd2",
X"3f83e080",
X"0856807d",
X"34838139",
X"933d841c",
X"08705859",
X"5f8a55a0",
X"76708105",
X"5834ff15",
X"5574ff2e",
X"098106ef",
X"3880705a",
X"5c887f08",
X"5f5a7b81",
X"1d7081ff",
X"06601370",
X"3370af32",
X"7030a073",
X"27718025",
X"07515152",
X"5b535e57",
X"557480e7",
X"3876ae2e",
X"09810683",
X"38815578",
X"7a277507",
X"5574802e",
X"9f387988",
X"32703078",
X"ae327030",
X"7073079f",
X"2a535157",
X"515675bb",
X"3888598b",
X"5affab39",
X"76982b55",
X"74802587",
X"3880f5c4",
X"173357ff",
X"9f175574",
X"99268938",
X"e0177081",
X"ff065855",
X"78811a70",
X"81ff0672",
X"1b535b57",
X"55767534",
X"fef8397b",
X"1e7f0c80",
X"5576a026",
X"83388155",
X"748b1934",
X"7a51fc82",
X"3f83e080",
X"0880f538",
X"a0547a22",
X"70852b83",
X"e0065455",
X"901b0852",
X"7c51a493",
X"3f83e080",
X"085783e0",
X"80088181",
X"387c3355",
X"74802e80",
X"f4388b1d",
X"3370832a",
X"70810651",
X"565674b4",
X"388b7d84",
X"1d0883e0",
X"8008595b",
X"5b58ff18",
X"5877ff2e",
X"9a387970",
X"81055b33",
X"79708105",
X"5b337171",
X"31525656",
X"75802ee2",
X"38863975",
X"802e9638",
X"7a51fbe5",
X"3fff8639",
X"83e08008",
X"5683e080",
X"08b63883",
X"39765684",
X"1b088b11",
X"33515574",
X"a7388b1d",
X"3370842a",
X"70810651",
X"56567489",
X"38835694",
X"39815690",
X"397c51fa",
X"943f83e0",
X"8008881c",
X"0cfd8139",
X"7583e080",
X"0c903d0d",
X"04f83d0d",
X"7a7c5957",
X"825483fe",
X"53775276",
X"51a2d83f",
X"835683e0",
X"800880ec",
X"38811733",
X"77337188",
X"2b075656",
X"82567482",
X"d4d52e09",
X"810680d4",
X"387554b6",
X"53775276",
X"51a2ac3f",
X"83e08008",
X"98388117",
X"33773371",
X"882b0783",
X"e0800852",
X"56567481",
X"82c62eac",
X"38825480",
X"d2537752",
X"7651a283",
X"3f83e080",
X"08983881",
X"17337733",
X"71882b07",
X"83e08008",
X"52565674",
X"8182c62e",
X"83388156",
X"7583e080",
X"0c8a3d0d",
X"04eb3d0d",
X"675a800b",
X"83e0900c",
X"a1a53f83",
X"e0800881",
X"06558256",
X"7483ef38",
X"7475538f",
X"3d705357",
X"59feca3f",
X"83e08008",
X"81ff0657",
X"76812e09",
X"810680d4",
X"38905483",
X"be537452",
X"7551a197",
X"3f83e080",
X"0880c938",
X"8f3d3355",
X"74802e80",
X"c93802bf",
X"05330284",
X"05be0533",
X"71982b71",
X"902b0702",
X"8c05bd05",
X"3370882b",
X"7207953d",
X"33710770",
X"587b575e",
X"525e5759",
X"57fdee3f",
X"83e08008",
X"81ff0657",
X"76832e09",
X"81068638",
X"815682f2",
X"3976802e",
X"86388656",
X"82e839a4",
X"548d5378",
X"527551a0",
X"ae3f8156",
X"83e08008",
X"82d43802",
X"be053302",
X"8405bd05",
X"3371882b",
X"07595d77",
X"ab380280",
X"ce053302",
X"840580cd",
X"05337198",
X"2b71902b",
X"07973d33",
X"70882b72",
X"07029405",
X"80cb0533",
X"71075452",
X"5e575956",
X"02b70533",
X"78712902",
X"8805b605",
X"33028c05",
X"b5053371",
X"882b0770",
X"1d707f8c",
X"050c5f59",
X"57595d8e",
X"3d33821b",
X"3402b905",
X"33903d33",
X"71882b07",
X"5a5c7884",
X"1b2302bb",
X"05330284",
X"05ba0533",
X"71882b07",
X"565c74ab",
X"380280ca",
X"05330284",
X"0580c905",
X"3371982b",
X"71902b07",
X"963d3370",
X"882b7207",
X"02940580",
X"c7053371",
X"07515253",
X"575e5c74",
X"76317831",
X"79842a90",
X"3d335471",
X"71315356",
X"5680d38a",
X"3f83e080",
X"08820570",
X"881c0c83",
X"e08008e0",
X"8a055656",
X"7483dffe",
X"26833882",
X"5783fff6",
X"76278538",
X"83578939",
X"86567680",
X"2e80db38",
X"767a3476",
X"832e0981",
X"06b03802",
X"80d60533",
X"02840580",
X"d5053371",
X"982b7190",
X"2b07993d",
X"3370882b",
X"72070294",
X"0580d305",
X"3371077f",
X"90050c52",
X"5e575856",
X"8639771b",
X"901b0c84",
X"1a228c1b",
X"08197184",
X"2a05941c",
X"0c5d800b",
X"811b3479",
X"83e0900c",
X"80567583",
X"e0800c97",
X"3d0d04e9",
X"3d0d83e0",
X"90085685",
X"5475802e",
X"81823880",
X"0b811734",
X"993de011",
X"466a548a",
X"3d705458",
X"ec0551f6",
X"e53f83e0",
X"80085483",
X"e0800880",
X"df38893d",
X"33547380",
X"2e913802",
X"ab053370",
X"842a8106",
X"51557480",
X"2e863883",
X"5480c139",
X"7651f489",
X"3f83e080",
X"08a0170c",
X"02bf0533",
X"028405be",
X"05337198",
X"2b71902b",
X"07028c05",
X"bd053370",
X"882b7207",
X"953d3371",
X"079c1c0c",
X"5278981b",
X"0c535659",
X"57810b81",
X"17347454",
X"7383e080",
X"0c993d0d",
X"04f53d0d",
X"7d7f6172",
X"83e09008",
X"5a5d5d59",
X"5c807b0c",
X"85577580",
X"2e81e038",
X"81163381",
X"06558457",
X"74802e81",
X"d2389139",
X"74811734",
X"8639800b",
X"81173481",
X"5781c039",
X"9c160898",
X"17083155",
X"74782783",
X"38745877",
X"802e81a9",
X"38981608",
X"7083ff06",
X"56577480",
X"cf388216",
X"33ff0577",
X"892a0670",
X"81ff065a",
X"5578a038",
X"768738a0",
X"1608558d",
X"39a41608",
X"51f0e93f",
X"83e08008",
X"55817527",
X"ffa83874",
X"a4170ca4",
X"160851f2",
X"833f83e0",
X"80085583",
X"e0800880",
X"2eff8938",
X"83e08008",
X"19a8170c",
X"98160883",
X"ff068480",
X"71315155",
X"77752783",
X"38775574",
X"83ffff06",
X"54981608",
X"83ff0653",
X"a8160852",
X"79577b83",
X"387b5776",
X"519ad43f",
X"83e08008",
X"fed03898",
X"16081598",
X"170c741a",
X"7876317c",
X"08177d0c",
X"595afed3",
X"39805776",
X"83e0800c",
X"8d3d0d04",
X"fa3d0d78",
X"83e09008",
X"55568555",
X"73802e81",
X"e3388114",
X"33810653",
X"84557280",
X"2e81d538",
X"9c140853",
X"72762783",
X"38725698",
X"14085780",
X"0b98150c",
X"75802e81",
X"b9388214",
X"3370892b",
X"56537680",
X"2eb73874",
X"52ff1651",
X"80ce8b3f",
X"83e08008",
X"ff187654",
X"70535853",
X"80cdfb3f",
X"83e08008",
X"73269638",
X"74307078",
X"06709817",
X"0c777131",
X"a4170852",
X"58515389",
X"39a01408",
X"70a4160c",
X"53747627",
X"b9387251",
X"eed63f83",
X"e0800853",
X"810b83e0",
X"8008278b",
X"38881408",
X"83e08008",
X"26883880",
X"0b811534",
X"b03983e0",
X"8008a415",
X"0c981408",
X"1598150c",
X"75753156",
X"c4399814",
X"08167098",
X"160c7352",
X"56efc53f",
X"83e08008",
X"8c3883e0",
X"80088115",
X"34815594",
X"39821433",
X"ff057689",
X"2a0683e0",
X"800805a8",
X"150c8055",
X"7483e080",
X"0c883d0d",
X"04ef3d0d",
X"63568555",
X"83e09008",
X"802e80d2",
X"38933df4",
X"0584170c",
X"6453883d",
X"70537652",
X"57f1cf3f",
X"83e08008",
X"5583e080",
X"08b43888",
X"3d335473",
X"802ea138",
X"02a70533",
X"70842a70",
X"81065155",
X"55835573",
X"802e9738",
X"7651eef5",
X"3f83e080",
X"0888170c",
X"7551efa6",
X"3f83e080",
X"08557483",
X"e0800c93",
X"3d0d04e4",
X"3d0d6ea1",
X"3d08405e",
X"855683e0",
X"9008802e",
X"8485389e",
X"3df40584",
X"1f0c7e98",
X"387d51ee",
X"f53f83e0",
X"80085683",
X"ee398141",
X"81f63983",
X"4181f139",
X"933d7f96",
X"05415980",
X"7f829505",
X"5e567560",
X"81ff0534",
X"8341901e",
X"08762e81",
X"d338a054",
X"7d227085",
X"2b83e006",
X"5458901e",
X"08527851",
X"96dd3f83",
X"e0800841",
X"83e08008",
X"ffb83878",
X"335c7b80",
X"2effb438",
X"8b193370",
X"bf067181",
X"06524355",
X"74802e80",
X"de387b81",
X"bf065574",
X"8f2480d3",
X"389a1933",
X"557480cb",
X"38f31d70",
X"585d8156",
X"758b2e09",
X"81068538",
X"8e568b39",
X"759a2e09",
X"81068338",
X"9c567519",
X"70708105",
X"52337133",
X"811a821a",
X"5f5b525b",
X"55748638",
X"79773485",
X"3980df77",
X"34777b57",
X"577aa02e",
X"098106c0",
X"3881567b",
X"81e53270",
X"30709f2a",
X"5151557b",
X"ae2e9338",
X"74802e8e",
X"3861832a",
X"70810651",
X"5574802e",
X"97387d51",
X"eddf3f83",
X"e0800841",
X"83e08008",
X"8738901e",
X"08feaf38",
X"80603475",
X"802e8838",
X"7c527f51",
X"8e833f60",
X"802e8638",
X"800b901f",
X"0c605660",
X"832e8538",
X"6081d038",
X"891f5790",
X"1e08802e",
X"81a83880",
X"56751970",
X"33515574",
X"a02ea038",
X"74852e09",
X"81068438",
X"81e55574",
X"77708105",
X"59348116",
X"7081ff06",
X"57558776",
X"27d73888",
X"19335574",
X"a02ea938",
X"ae777081",
X"05593488",
X"56751970",
X"33515574",
X"a02e9538",
X"74777081",
X"05593481",
X"167081ff",
X"0657558a",
X"7627e238",
X"8b19337f",
X"8805349f",
X"19339e1a",
X"3371982b",
X"71902b07",
X"9d1c3370",
X"882b7207",
X"9c1e3371",
X"07640c52",
X"991d3398",
X"1e337188",
X"2b075351",
X"53575956",
X"747f8405",
X"23971933",
X"961a3371",
X"882b0756",
X"56747f86",
X"05238077",
X"347d51eb",
X"f03f83e0",
X"80088332",
X"70307072",
X"079f2c83",
X"e0800806",
X"52565696",
X"1f335574",
X"8a38891f",
X"52961f51",
X"8c8f3f75",
X"83e0800c",
X"9e3d0d04",
X"f43d0d7e",
X"8f3dec11",
X"56565890",
X"53f01552",
X"7751e0d2",
X"3f83e080",
X"0880d738",
X"78902e09",
X"810680ce",
X"3802ab05",
X"3380fb80",
X"0b80fb80",
X"33575856",
X"8c397476",
X"2e8a3884",
X"17703356",
X"5774f338",
X"76337057",
X"5574802e",
X"ad388217",
X"22708a2b",
X"903dec05",
X"56705556",
X"56848880",
X"80527751",
X"e0803f83",
X"e0800886",
X"3878752e",
X"85388056",
X"85398117",
X"33567583",
X"e0800c8e",
X"3d0d04fc",
X"3d0d7670",
X"52558b95",
X"3f83e080",
X"0815ff05",
X"5473752e",
X"8e387333",
X"5372ae2e",
X"8638ff14",
X"54ef3977",
X"52811451",
X"8aad3f83",
X"e0800830",
X"7083e080",
X"08078025",
X"83e0800c",
X"53863d0d",
X"04fc3d0d",
X"76705255",
X"e6ed3f83",
X"e0800854",
X"815383e0",
X"800880c1",
X"387451e6",
X"b03f83e0",
X"800880f8",
X"845383e0",
X"80085253",
X"ff913f83",
X"e08008a1",
X"3880f888",
X"527251ff",
X"823f83e0",
X"80089238",
X"80f88c52",
X"7251fef3",
X"3f83e080",
X"08802e83",
X"38815473",
X"537283e0",
X"800c863d",
X"0d04fd3d",
X"0d757052",
X"54e68c3f",
X"815383e0",
X"80089838",
X"7351e5d5",
X"3f83e388",
X"085283e0",
X"800851fe",
X"ba3f83e0",
X"80085372",
X"83e0800c",
X"853d0d04",
X"df3d0da4",
X"3d087052",
X"5edbfa3f",
X"83e08008",
X"33953d56",
X"54739638",
X"80febc52",
X"7451898d",
X"3f9a397d",
X"527851de",
X"fb3f84d0",
X"397d51db",
X"e03f83e0",
X"80085274",
X"51db903f",
X"80438042",
X"80418040",
X"83e39008",
X"52943d70",
X"525de1e3",
X"3f83e080",
X"0859800b",
X"83e08008",
X"555b83e0",
X"80087b2e",
X"9438811b",
X"74525be4",
X"e53f83e0",
X"80085483",
X"e08008ee",
X"38805aff",
X"5f790970",
X"9f2c7b06",
X"5b547a7a",
X"248438ff",
X"1b5af61a",
X"7009709f",
X"2c72067b",
X"ff125a5a",
X"52555580",
X"75259538",
X"7651e4aa",
X"3f83e080",
X"0876ff18",
X"58555773",
X"8024ed38",
X"747f2e86",
X"38a1b53f",
X"745f78ff",
X"1b70585d",
X"58807a25",
X"95387751",
X"e4803f83",
X"e0800876",
X"ff185855",
X"58738024",
X"ed38800b",
X"83e7c00c",
X"800b83e7",
X"e40c80f8",
X"90518d8c",
X"3f81800b",
X"83e7e40c",
X"80f89851",
X"8cfe3fa8",
X"0b83e7c0",
X"0c76802e",
X"80e43883",
X"e7c00877",
X"79327030",
X"70720780",
X"2570872b",
X"83e7e40c",
X"51567853",
X"5656e3b7",
X"3f83e080",
X"08802e88",
X"3880f8a0",
X"518cc53f",
X"7651e2f9",
X"3f83e080",
X"085280f9",
X"c0518cb4",
X"3f7651e3",
X"813f83e0",
X"800883e7",
X"c0085557",
X"75742586",
X"38a81656",
X"f7397583",
X"e7c00c86",
X"f07624ff",
X"98388798",
X"0b83e7c0",
X"0c77802e",
X"b1387751",
X"e2b73f83",
X"e0800878",
X"5255e2d7",
X"3f80f8a8",
X"5483e080",
X"088d3887",
X"39807634",
X"81d03980",
X"f8a45474",
X"53735280",
X"f7f8518b",
X"d33f8054",
X"80f88051",
X"8bca3f81",
X"145473a8",
X"2e098106",
X"ef38868d",
X"a0519da8",
X"3f805290",
X"3d705257",
X"80c3ef3f",
X"83527651",
X"80c3e73f",
X"62818f38",
X"61802e80",
X"fb387b54",
X"73ff2e96",
X"3878802e",
X"818a3878",
X"51e1db3f",
X"83e08008",
X"ff155559",
X"e7397880",
X"2e80f538",
X"7851e1d7",
X"3f83e080",
X"08802efc",
X"8e387851",
X"e19f3f83",
X"e0800852",
X"80f7f451",
X"83e03f83",
X"e08008a3",
X"387c5185",
X"983f83e0",
X"80085574",
X"ff165654",
X"807425ae",
X"38741d70",
X"33555673",
X"af2efecd",
X"38e93978",
X"51e0e03f",
X"83e08008",
X"527c5184",
X"d03f8f39",
X"7f882960",
X"10057a05",
X"61055afc",
X"90396280",
X"2efbd138",
X"80527651",
X"80c2c73f",
X"a33d0d04",
X"803d0d90",
X"88b83370",
X"81ff0670",
X"842a8132",
X"70810651",
X"51515170",
X"802e8d38",
X"a80b9088",
X"b834b80b",
X"9088b834",
X"7083e080",
X"0c823d0d",
X"04803d0d",
X"9088b833",
X"7081ff06",
X"70852a81",
X"32708106",
X"51515151",
X"70802e8d",
X"38980b90",
X"88b834b8",
X"0b9088b8",
X"347083e0",
X"800c823d",
X"0d04930b",
X"9088bc34",
X"ff0b9088",
X"a83404ff",
X"3d0d028f",
X"05335280",
X"0b9088bc",
X"348a519a",
X"ef3fdf3f",
X"80f80b90",
X"88a03480",
X"0b908888",
X"34fa1252",
X"71908880",
X"34800b90",
X"88983471",
X"90889034",
X"9088b852",
X"807234b8",
X"7234833d",
X"0d04803d",
X"0d028b05",
X"33517090",
X"88b434fe",
X"bf3f83e0",
X"8008802e",
X"f638823d",
X"0d04803d",
X"0d8439a6",
X"ac3ffed9",
X"3f83e080",
X"08802ef3",
X"389088b4",
X"337081ff",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0da30b90",
X"88bc34ff",
X"0b9088a8",
X"349088b8",
X"51a87134",
X"b8713482",
X"3d0d0480",
X"3d0d9088",
X"bc337098",
X"2b708025",
X"83e0800c",
X"5151823d",
X"0d04803d",
X"0d9088b8",
X"337081ff",
X"0670832a",
X"81327081",
X"06515151",
X"5170802e",
X"e838b00b",
X"9088b834",
X"b80b9088",
X"b834823d",
X"0d04803d",
X"0d9080ac",
X"08810683",
X"e0800c82",
X"3d0d04fd",
X"3d0d7577",
X"54548073",
X"25943873",
X"70810555",
X"335280f8",
X"ac518784",
X"3fff1353",
X"e939853d",
X"0d04fd3d",
X"0d757753",
X"54733351",
X"70893871",
X"33517080",
X"2ea13873",
X"33723352",
X"53727127",
X"8538ff51",
X"94397073",
X"27853881",
X"518b3981",
X"14811353",
X"54d33980",
X"517083e0",
X"800c853d",
X"0d04fd3d",
X"0d757754",
X"54723370",
X"81ff0652",
X"5270802e",
X"a3387181",
X"ff068114",
X"ffbf1253",
X"54527099",
X"268938a0",
X"127081ff",
X"06535171",
X"74708105",
X"5634d239",
X"80743485",
X"3d0d04ff",
X"bd3d0d80",
X"c63d0852",
X"a53d7052",
X"54ffb33f",
X"80c73d08",
X"52853d70",
X"5253ffa6",
X"3f725273",
X"51fedf3f",
X"80c53d0d",
X"04fe3d0d",
X"74765353",
X"71708105",
X"53335170",
X"73708105",
X"553470f0",
X"38843d0d",
X"04fe3d0d",
X"74528072",
X"33525370",
X"732e8d38",
X"81128114",
X"71335354",
X"5270f538",
X"7283e080",
X"0c843d0d",
X"04f63d0d",
X"7c7e6062",
X"5a5d5b56",
X"80598155",
X"8539747a",
X"29557452",
X"7551bae2",
X"3f83e080",
X"087a27ee",
X"3874802e",
X"80dd3874",
X"527551ba",
X"cd3f83e0",
X"80087553",
X"765254ba",
X"d13f83e0",
X"80087a53",
X"755256ba",
X"b53f83e0",
X"80087930",
X"707b079f",
X"2a707780",
X"24075151",
X"54557287",
X"3883e080",
X"08c53876",
X"8118b016",
X"55585889",
X"74258b38",
X"b714537a",
X"853880d7",
X"14537278",
X"34811959",
X"ff9f3980",
X"77348c3d",
X"0d04f73d",
X"0d7b7d7f",
X"62029005",
X"bb053357",
X"59565a5a",
X"b0587283",
X"38a05875",
X"70708105",
X"52337159",
X"54559039",
X"8074258e",
X"38ff1477",
X"70810559",
X"33545472",
X"ef3873ff",
X"15555380",
X"73258938",
X"77527951",
X"782def39",
X"75337557",
X"5372802e",
X"90387252",
X"7951782d",
X"75708105",
X"573353ed",
X"398b3d0d",
X"04ee3d0d",
X"64666969",
X"70708105",
X"52335b4a",
X"5c5e5e76",
X"802e82f9",
X"3876a52e",
X"09810682",
X"e0388070",
X"41677070",
X"81055233",
X"714a5957",
X"5f76b02e",
X"0981068c",
X"38757081",
X"05573376",
X"4857815f",
X"d0175675",
X"892680da",
X"3876675c",
X"59805c93",
X"39778a24",
X"80c3387b",
X"8a29187b",
X"7081055d",
X"335a5cd0",
X"197081ff",
X"06585889",
X"7727a438",
X"ff9f1970",
X"81ff06ff",
X"a91b5a51",
X"56857627",
X"9238ffbf",
X"197081ff",
X"06515675",
X"85268a38",
X"c9195877",
X"8025ffb9",
X"387a477b",
X"407881ff",
X"06577680",
X"e42e80e5",
X"387680e4",
X"24a73876",
X"80d82e81",
X"86387680",
X"d8249038",
X"76802e81",
X"cc3876a5",
X"2e81b638",
X"81b93976",
X"80e32e81",
X"8c3881af",
X"397680f5",
X"2e9b3876",
X"80f5248b",
X"387680f3",
X"2e818138",
X"81993976",
X"80f82e80",
X"ca38818f",
X"39913d70",
X"55578053",
X"8a527984",
X"1b710853",
X"5b56fc81",
X"3f7655ab",
X"3979841b",
X"7108943d",
X"705b5b52",
X"5b567580",
X"258c3875",
X"3056ad78",
X"340280c1",
X"05577654",
X"80538a52",
X"7551fbd5",
X"3f77557e",
X"54b83991",
X"3d705577",
X"80d83270",
X"30708025",
X"56515856",
X"90527984",
X"1b710853",
X"5b57fbb1",
X"3f7555db",
X"3979841b",
X"83123354",
X"5b569839",
X"79841b71",
X"08575b56",
X"80547f53",
X"7c527d51",
X"fc9c3f87",
X"3976527d",
X"517c2d66",
X"70335881",
X"0547fd83",
X"39943d0d",
X"047283e0",
X"940c7183",
X"e0980c04",
X"fb3d0d88",
X"3d707084",
X"05520857",
X"54755383",
X"e0940852",
X"83e09808",
X"51fcc63f",
X"873d0d04",
X"ff3d0d73",
X"70085351",
X"02930533",
X"72347008",
X"8105710c",
X"833d0d04",
X"fc3d0d87",
X"3d881155",
X"7854bdb8",
X"5351fc99",
X"3f805287",
X"3d51d13f",
X"863d0d04",
X"fc3d0d76",
X"557483e3",
X"9c082eaf",
X"38805374",
X"5187c13f",
X"83e08008",
X"81ff06ff",
X"147081ff",
X"06723070",
X"9f2a5152",
X"55535472",
X"802e8438",
X"71dd3873",
X"fe387483",
X"e39c0c86",
X"3d0d04ff",
X"3d0dff0b",
X"83e39c0c",
X"84a53f81",
X"5187853f",
X"83e08008",
X"81ff0652",
X"71ee3881",
X"d33f7183",
X"e0800c83",
X"3d0d04fc",
X"3d0d7602",
X"8405a205",
X"22028805",
X"a605227a",
X"54555555",
X"ff823f72",
X"802ea038",
X"83e3b014",
X"33757081",
X"05573481",
X"147083ff",
X"ff06ff15",
X"7083ffff",
X"06565255",
X"52dd3980",
X"0b83e080",
X"0c863d0d",
X"04fc3d0d",
X"76787a11",
X"56535580",
X"5371742e",
X"93387215",
X"51703383",
X"e3b01334",
X"81128114",
X"5452ea39",
X"800b83e0",
X"800c863d",
X"0d04fd3d",
X"0d905483",
X"e39c0851",
X"86f43f83",
X"e0800881",
X"ff06ff15",
X"71307130",
X"7073079f",
X"2a729f2a",
X"06525552",
X"555372db",
X"38853d0d",
X"04803d0d",
X"83e3a808",
X"1083e3a0",
X"08079080",
X"a80c823d",
X"0d04800b",
X"83e3a80c",
X"e43f0481",
X"0b83e3a8",
X"0cdb3f04",
X"ed3f0471",
X"83e3a40c",
X"04803d0d",
X"8051f43f",
X"810b83e3",
X"a80c810b",
X"83e3a00c",
X"ffbb3f82",
X"3d0d0480",
X"3d0d7230",
X"70740780",
X"2583e3a0",
X"0c51ffa5",
X"3f823d0d",
X"04803d0d",
X"028b0533",
X"9080a40c",
X"9080a808",
X"70810651",
X"5170f538",
X"9080a408",
X"7081ff06",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"81ff51d1",
X"3f83e080",
X"0881ff06",
X"83e0800c",
X"823d0d04",
X"803d0d73",
X"902b7307",
X"9080b40c",
X"823d0d04",
X"04fb3d0d",
X"78028405",
X"9f053370",
X"982b5557",
X"55728025",
X"9b387580",
X"ff065680",
X"5280f751",
X"e03f83e0",
X"800881ff",
X"06547381",
X"2680ff38",
X"8051fee7",
X"3fffa23f",
X"8151fedf",
X"3fff9a3f",
X"7551feed",
X"3f74982a",
X"51fee63f",
X"74902a70",
X"81ff0652",
X"53feda3f",
X"74882a70",
X"81ff0652",
X"53fece3f",
X"7481ff06",
X"51fec63f",
X"81557580",
X"c02e0981",
X"06863881",
X"95558d39",
X"7580c82e",
X"09810684",
X"38818755",
X"7451fea5",
X"3f8a55fe",
X"c83f83e0",
X"800881ff",
X"0670982b",
X"54547280",
X"258c38ff",
X"157081ff",
X"06565374",
X"e2387383",
X"e0800c87",
X"3d0d04fa",
X"3d0dfdc5",
X"3f8051fd",
X"da3f8a54",
X"fe933fff",
X"147081ff",
X"06555373",
X"f3387374",
X"535580c0",
X"51fea63f",
X"83e08008",
X"81ff0654",
X"73812e09",
X"8106829f",
X"3883aa52",
X"80c851fe",
X"8c3f83e0",
X"800881ff",
X"06537281",
X"2e098106",
X"81a83874",
X"54873d74",
X"115456fd",
X"c83f83e0",
X"80087334",
X"81147081",
X"ff065553",
X"837427e5",
X"38029a05",
X"33537281",
X"2e098106",
X"81d93802",
X"9b053353",
X"80ce9054",
X"7281aa2e",
X"8d3881c7",
X"3980e451",
X"8b9a3fff",
X"14547380",
X"2e81b838",
X"820a5281",
X"e951fda5",
X"3f83e080",
X"0881ff06",
X"5372de38",
X"725280fa",
X"51fd923f",
X"83e08008",
X"81ff0653",
X"72819038",
X"72547316",
X"53fcd63f",
X"83e08008",
X"73348114",
X"7081ff06",
X"55538374",
X"27e83887",
X"3d337086",
X"2a708106",
X"5154548c",
X"557280e3",
X"38845580",
X"de397452",
X"81e951fc",
X"cc3f83e0",
X"800881ff",
X"06538255",
X"81e95681",
X"73278638",
X"735580c1",
X"5680ce90",
X"548a3980",
X"e4518a8c",
X"3fff1454",
X"73802ea9",
X"38805275",
X"51fc9a3f",
X"83e08008",
X"81ff0653",
X"72e13884",
X"805280d0",
X"51fc863f",
X"83e08008",
X"81ff0653",
X"72802e83",
X"38805574",
X"83e3ac34",
X"8051fb87",
X"3ffbc23f",
X"883d0d04",
X"fb3d0d77",
X"54800b83",
X"e3ac3370",
X"832a7081",
X"06515557",
X"5572752e",
X"09810685",
X"3873892b",
X"54735280",
X"d151fbbd",
X"3f83e080",
X"0881ff06",
X"5372bd38",
X"82b8c054",
X"fb833f83",
X"e0800881",
X"ff065372",
X"81ff2e09",
X"81068938",
X"ff145473",
X"e7389f39",
X"7281fe2e",
X"09810696",
X"3883e7b0",
X"5283e3b0",
X"51faed3f",
X"fad33ffa",
X"d03f8339",
X"81558051",
X"fa893ffa",
X"c43f7481",
X"ff0683e0",
X"800c873d",
X"0d04fb3d",
X"0d7783e3",
X"b0565481",
X"51f9ec3f",
X"83e3ac33",
X"70832a70",
X"81065154",
X"56728538",
X"73892b54",
X"735280d8",
X"51fab63f",
X"83e08008",
X"81ff0653",
X"7280e438",
X"81ff51f9",
X"d43f81fe",
X"51f9ce3f",
X"84805374",
X"70810556",
X"3351f9c1",
X"3fff1370",
X"83ffff06",
X"515372eb",
X"387251f9",
X"b03f7251",
X"f9ab3ff9",
X"d03f83e0",
X"80089f06",
X"53a78854",
X"72852e8c",
X"38993980",
X"e45187c4",
X"3fff1454",
X"f9b33f83",
X"e0800881",
X"ff2e8438",
X"73e93880",
X"51f8e43f",
X"f99f3f80",
X"0b83e080",
X"0c873d0d",
X"047183e7",
X"b40c8880",
X"800b83e7",
X"b00c8480",
X"800b83e7",
X"b80c04fd",
X"3d0d7770",
X"17557705",
X"ff1a5353",
X"71ff2e94",
X"38737081",
X"05553351",
X"70737081",
X"055534ff",
X"1252e939",
X"853d0d04",
X"fb3d0d87",
X"a6810b83",
X"e7b40856",
X"56753383",
X"a6801634",
X"a05483a0",
X"805383e7",
X"b4085283",
X"e7b00851",
X"ffb13fa0",
X"5483a480",
X"5383e7b4",
X"085283e7",
X"b00851ff",
X"9e3f9054",
X"83a88053",
X"83e7b408",
X"5283e7b0",
X"0851ff8b",
X"3fa05380",
X"5283e7b8",
X"0883a080",
X"05518695",
X"3fa05380",
X"5283e7b8",
X"0883a480",
X"05518685",
X"3f905380",
X"5283e7b8",
X"0883a880",
X"055185f5",
X"3fff7634",
X"83a08054",
X"805383e7",
X"b4085283",
X"e7b80851",
X"fec53f80",
X"d0805483",
X"b0805383",
X"e7b40852",
X"83e7b808",
X"51feb03f",
X"87ba3fa2",
X"54805383",
X"e7b8088c",
X"80055280",
X"fbf451fe",
X"9a3f860b",
X"87a88334",
X"800b87a8",
X"8234800b",
X"87a09a34",
X"af0b87a0",
X"9634bf0b",
X"87a09734",
X"800b87a0",
X"98349f0b",
X"87a09934",
X"800b87a0",
X"9b34e00b",
X"87a88934",
X"a20b87a8",
X"8034830b",
X"87a48f34",
X"820b87a8",
X"8134873d",
X"0d04fc3d",
X"0d83a080",
X"54805383",
X"e7b80852",
X"83e7b408",
X"51fdb83f",
X"80d08054",
X"83b08053",
X"83e7b808",
X"5283e7b4",
X"0851fda3",
X"3fa05483",
X"a0805383",
X"e7b80852",
X"83e7b408",
X"51fd903f",
X"a05483a4",
X"805383e7",
X"b8085283",
X"e7b40851",
X"fcfd3f90",
X"5483a880",
X"5383e7b8",
X"085283e7",
X"b40851fc",
X"ea3f83e7",
X"b4085583",
X"a6801533",
X"87a68134",
X"863d0d04",
X"fa3d0d78",
X"705255c1",
X"e23f83ff",
X"ff0b83e0",
X"800825a9",
X"387451c1",
X"e33f83e0",
X"80089e38",
X"83e08008",
X"57883dfc",
X"05548480",
X"805383e7",
X"b4085274",
X"51ffbf9c",
X"3fffbee2",
X"3f883d0d",
X"04fa3d0d",
X"78705255",
X"c1a13f83",
X"ffff0b83",
X"e0800825",
X"96388057",
X"883dfc05",
X"54848080",
X"5383e7b4",
X"08527451",
X"c0943f88",
X"3d0d0480",
X"3d0d9080",
X"90088106",
X"83e0800c",
X"823d0d04",
X"ff3d0d90",
X"80907008",
X"70fe0676",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70812c81",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870fd",
X"06761007",
X"720c5252",
X"833d0d04",
X"803d0d90",
X"80900870",
X"822cbf06",
X"83e0800c",
X"51823d0d",
X"04ff3d0d",
X"90809070",
X"0870fe83",
X"0676822b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70882c87",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870f1",
X"ff067688",
X"2b07720c",
X"5252833d",
X"0d04803d",
X"0d908090",
X"0870912c",
X"bf0683e0",
X"800c5182",
X"3d0d04ff",
X"3d0d9080",
X"90700870",
X"fc87ffff",
X"0676912b",
X"07720c52",
X"52833d0d",
X"04803d0d",
X"90809008",
X"70992c81",
X"0683e080",
X"0c51823d",
X"0d04ff3d",
X"0d908090",
X"700870ff",
X"bf0a0676",
X"992b0772",
X"0c525283",
X"3d0d0480",
X"3d0d9080",
X"80087088",
X"2c810683",
X"e0800c51",
X"823d0d04",
X"803d0d90",
X"80800870",
X"892c8106",
X"83e0800c",
X"51823d0d",
X"04803d0d",
X"90808008",
X"708a2c81",
X"0683e080",
X"0c51823d",
X"0d04803d",
X"0d908080",
X"08708b2c",
X"810683e0",
X"800c5182",
X"3d0d0480",
X"3d0d9080",
X"8008708c",
X"2cbf0683",
X"e0800c51",
X"823d0d04",
X"fe3d0d74",
X"81e62987",
X"2a9080a0",
X"0c843d0d",
X"04fe3d0d",
X"7575ff19",
X"53535370",
X"ff2e8d38",
X"72727081",
X"055434ff",
X"1151f039",
X"843d0d04",
X"fe3d0d75",
X"75ff1953",
X"535370ff",
X"2e8d3872",
X"72708405",
X"540cff11",
X"51f03984",
X"3d0d04fe",
X"3d0d8480",
X"80538052",
X"88800a51",
X"ffb33f81",
X"80805380",
X"5282800a",
X"51c63f84",
X"3d0d0480",
X"3d0d8151",
X"fcaa3f72",
X"802e9038",
X"8051fdfe",
X"3fcd3f83",
X"e7bc3351",
X"fdf43f81",
X"51fcbb3f",
X"8051fcb6",
X"3f8051fc",
X"873f823d",
X"0d04fd3d",
X"0d755280",
X"5480ff72",
X"25883881",
X"0bff8013",
X"5354ffbf",
X"12517099",
X"268638e0",
X"1252b039",
X"ff9f1251",
X"997127a7",
X"38d012e0",
X"13545170",
X"89268538",
X"72529839",
X"728f2685",
X"3872528f",
X"3971ba2e",
X"09810685",
X"389a5283",
X"39805273",
X"802e8538",
X"81801252",
X"7181ff06",
X"83e0800c",
X"853d0d04",
X"803d0d84",
X"d8c05180",
X"71708105",
X"53347084",
X"e0c02e09",
X"8106f038",
X"823d0d04",
X"fe3d0d02",
X"97053351",
X"fef43f83",
X"e0800881",
X"ff0683e7",
X"c0085452",
X"8073249b",
X"3883e7e0",
X"08137283",
X"e7e40807",
X"53537173",
X"3483e7c0",
X"08810583",
X"e7c00c84",
X"3d0d04fa",
X"3d0d8280",
X"0a1b5580",
X"57883dfc",
X"05547953",
X"74527851",
X"ffbaab3f",
X"883d0d04",
X"fe3d0d83",
X"e7d80852",
X"7451c18f",
X"3f83e080",
X"088c3876",
X"53755283",
X"e7d80851",
X"c63f843d",
X"0d04fe3d",
X"0d83e7d8",
X"08537552",
X"7451ffbb",
X"cd3f83e0",
X"80088d38",
X"77537652",
X"83e7d808",
X"51ffa03f",
X"843d0d04",
X"fe3d0d83",
X"e7d80851",
X"ffbac03f",
X"83e08008",
X"8180802e",
X"09810687",
X"388f8080",
X"539b3983",
X"e7d80851",
X"ffbaa43f",
X"83e08008",
X"80d0802e",
X"09810692",
X"388fb080",
X"5383e080",
X"085283e7",
X"d80851fe",
X"d63f843d",
X"0d04803d",
X"0df9fe3f",
X"83e08008",
X"842980fc",
X"98057008",
X"83e0800c",
X"51823d0d",
X"04ed3d0d",
X"80448043",
X"80428041",
X"80705a5b",
X"fdce3f80",
X"0b83e7c0",
X"0c800b83",
X"e7e40c80",
X"f8f851e9",
X"c73f8180",
X"0b83e7e4",
X"0c80f8fc",
X"51e9b93f",
X"80d00b83",
X"e7c00c78",
X"30707a07",
X"80257087",
X"2b83e7e4",
X"0c5155f8",
X"ef3f83e0",
X"80085280",
X"f98451e9",
X"933f80f8",
X"0b83e7c0",
X"0c788132",
X"70307072",
X"07802570",
X"872b83e7",
X"e40c5156",
X"569df53f",
X"83e08008",
X"5280f994",
X"51e8e93f",
X"81a00b83",
X"e7c00c78",
X"82327030",
X"70720780",
X"2570872b",
X"83e7e40c",
X"515656fe",
X"c53f83e0",
X"80085280",
X"f9a451e8",
X"bf3f81c8",
X"0b83e7c0",
X"0c788332",
X"70307072",
X"07802570",
X"872b83e7",
X"e40c5156",
X"83e7d808",
X"5256ffb5",
X"a03f83e0",
X"80085280",
X"f9ac51e8",
X"8f3f8298",
X"0b83e7c0",
X"0c810b83",
X"e7c45b58",
X"83e7c008",
X"83197a32",
X"70307072",
X"07802570",
X"872b83e7",
X"e40c5157",
X"8e3d7055",
X"ff1b5457",
X"57579bb7",
X"3f797084",
X"055b0851",
X"ffb4d63f",
X"745483e0",
X"80085377",
X"5280f9b4",
X"51e7c13f",
X"a81783e7",
X"c00c8118",
X"5877852e",
X"098106ff",
X"af3883b8",
X"0b83e7c0",
X"0c788832",
X"70307072",
X"07802570",
X"872b83e7",
X"e40c5156",
X"56f7bb3f",
X"80f9c455",
X"83e08008",
X"802e8f38",
X"83e7d408",
X"51ffb481",
X"3f83e080",
X"08557452",
X"80f9cc51",
X"e6ee3f84",
X"880b83e7",
X"c00c7889",
X"32703070",
X"72078025",
X"70872b83",
X"e7e40c51",
X"5680f9d8",
X"5256e6cc",
X"3f84b00b",
X"83e7c00c",
X"788a3270",
X"30707207",
X"80257087",
X"2b83e7e4",
X"0c515680",
X"f9e45256",
X"e6aa3f85",
X"800b83e7",
X"c00c788b",
X"32703070",
X"72078025",
X"70872b83",
X"e7e40c51",
X"5680fa80",
X"5256e688",
X"3f868da0",
X"51f7f13f",
X"8052913d",
X"7052559e",
X"b93f8352",
X"74519eb2",
X"3f635574",
X"83e03861",
X"19597880",
X"25853874",
X"5990398b",
X"79258538",
X"8b598739",
X"788b2683",
X"bf387882",
X"2b5580f7",
X"c4150804",
X"f5923f83",
X"e0800861",
X"57557581",
X"2e098106",
X"893883e0",
X"80081055",
X"903975ff",
X"2e098106",
X"883883e0",
X"8008812c",
X"55907525",
X"85389055",
X"88397480",
X"24833881",
X"557451f4",
X"ec3f82f4",
X"3999f83f",
X"83e08008",
X"61055574",
X"80258538",
X"80558839",
X"87752583",
X"38875574",
X"518ddb3f",
X"82d239f4",
X"dc3f83e0",
X"80086105",
X"55748025",
X"85388055",
X"88398375",
X"25833883",
X"557451f4",
X"d53f82b0",
X"39608738",
X"62802e82",
X"a73883e3",
X"8c0883e3",
X"880cade6",
X"0b83e390",
X"0c83e7d8",
X"0851d5a0",
X"3ff9cd3f",
X"828a3960",
X"56807625",
X"9838ad85",
X"0b83e390",
X"0c83e7b4",
X"15700852",
X"55d5813f",
X"74085292",
X"39758025",
X"923883e7",
X"b4150851",
X"ffb1843f",
X"8052fc19",
X"51b83962",
X"802e81d0",
X"3883e7b4",
X"15700883",
X"e7c40872",
X"0c83e7c4",
X"0cfc1a70",
X"5351558c",
X"a83f83e0",
X"80085680",
X"518c9e3f",
X"83e08008",
X"52745188",
X"b73f7552",
X"805188b0",
X"3f819939",
X"60558075",
X"25b83883",
X"e3980883",
X"e3880cad",
X"e60b83e3",
X"900c83e7",
X"d40851d4",
X"8b3f83e7",
X"d40851d1",
X"ab3f83e0",
X"800881ff",
X"06705255",
X"f3b53f74",
X"802e80e0",
X"38815580",
X"e3397480",
X"2580d538",
X"83e7d408",
X"51ffaff3",
X"3f8051f3",
X"963f80c4",
X"3962802e",
X"bf3883e3",
X"940883e3",
X"880cade6",
X"0b83e390",
X"0c83e7dc",
X"0851d3b8",
X"3f78892e",
X"0981068b",
X"3883e7dc",
X"0851f0f9",
X"3f963978",
X"8a2e0981",
X"068e3883",
X"e7dc0851",
X"f0a63f84",
X"39628738",
X"7a802ef8",
X"af388055",
X"7483e080",
X"0c953d0d",
X"04fe3d0d",
X"f3813f83",
X"e0800880",
X"2e863880",
X"51818a39",
X"f3863f83",
X"e0800880",
X"fe38f3a6",
X"3f83e080",
X"08802eb9",
X"388151f0",
X"e33f8051",
X"f2bc3fec",
X"db3f800b",
X"83e7c00c",
X"f7d73f83",
X"e0800853",
X"ff0b83e7",
X"c00ceece",
X"3f7280cb",
X"3883e7bc",
X"3351f296",
X"3f7251f0",
X"b33f80c0",
X"39f2ce3f",
X"83e08008",
X"802eb538",
X"8151f0a0",
X"3f8051f1",
X"f93fec98",
X"3fad850b",
X"83e3900c",
X"83e7c408",
X"51d1f93f",
X"ff0b83e7",
X"c00cee8a",
X"3f83e7c4",
X"08528051",
X"85ea3f81",
X"51f3c03f",
X"843d0d04",
X"fc3d0d80",
X"0b83e7bc",
X"34848080",
X"52848a80",
X"8051ffb1",
X"eb3f83e0",
X"800880cd",
X"3889cf3f",
X"80feac51",
X"ffb6aa3f",
X"83e08008",
X"558e8080",
X"5480c080",
X"5380fa88",
X"5283e080",
X"0851f5a6",
X"3f83e7d8",
X"085380fa",
X"98527451",
X"ffb0f33f",
X"83e08008",
X"8438f5b4",
X"3f83e7bc",
X"3351f0ea",
X"3f8151f2",
X"d63f93ca",
X"3f8151f2",
X"ce3f8151",
X"fdeb3ffa",
X"3983e08c",
X"080283e0",
X"8c0cfb3d",
X"0d0280fa",
X"a40b83e3",
X"8c0c80fa",
X"a80b83e3",
X"840c80fa",
X"ac0b83e3",
X"980c80fa",
X"b00b83e3",
X"940c83e0",
X"8c08fc05",
X"0c800b83",
X"e7c40b83",
X"e08c08f8",
X"050c83e0",
X"8c08f405",
X"0cffafb8",
X"3f83e080",
X"088605fc",
X"0683e08c",
X"08f0050c",
X"0283e08c",
X"08f00508",
X"310d833d",
X"7083e08c",
X"08f80508",
X"70840583",
X"e08c08f8",
X"050c0c51",
X"ffac803f",
X"83e08c08",
X"f4050881",
X"0583e08c",
X"08f4050c",
X"83e08c08",
X"f4050887",
X"2e098106",
X"ffab3884",
X"84808051",
X"e9933fff",
X"0b83e7c0",
X"0c800b83",
X"e7e40c84",
X"d8c00b83",
X"e7e00c81",
X"51edb93f",
X"8151edde",
X"3f8051ed",
X"d93f8151",
X"edff3f82",
X"51eea73f",
X"8051eecf",
X"3f8051ee",
X"f93f80d1",
X"a8528051",
X"ddf73ffd",
X"a33f83e0",
X"8c08fc05",
X"080d800b",
X"83e0800c",
X"873d0d83",
X"e08c0c04",
X"803d0d81",
X"ff51800b",
X"83e7f412",
X"34ff1151",
X"70f43882",
X"3d0d04ff",
X"3d0d7370",
X"33535181",
X"11337134",
X"71811234",
X"833d0d04",
X"ff3d0d83",
X"ea9008a8",
X"2e098106",
X"8b3883ea",
X"a80883ea",
X"900c8739",
X"a80b83ea",
X"900c83ea",
X"90088605",
X"7081ff06",
X"5252d3ff",
X"3f833d0d",
X"04fb3d0d",
X"77795656",
X"80707155",
X"55527175",
X"25ac3872",
X"16703370",
X"147081ff",
X"06555151",
X"51717427",
X"89388112",
X"7081ff06",
X"53517181",
X"147083ff",
X"ff065552",
X"54747324",
X"d6387183",
X"e0800c87",
X"3d0d04fb",
X"3d0d7756",
X"8939fabd",
X"3f8351ee",
X"a73fd586",
X"3f83e080",
X"08802eee",
X"3883ea90",
X"08860570",
X"81ff0652",
X"53d38c3f",
X"810b9088",
X"d434fa95",
X"3f8351ed",
X"ff3f9088",
X"d4337081",
X"ff065553",
X"73802eea",
X"3873862a",
X"70810651",
X"5372ffbe",
X"3873982b",
X"53807324",
X"80de38d3",
X"f63f83e0",
X"80085583",
X"e0800880",
X"cf387416",
X"75822b54",
X"549088c0",
X"13337434",
X"81155574",
X"852e0981",
X"06e83875",
X"3383e7f4",
X"34811633",
X"83e7f534",
X"82163383",
X"e7f63483",
X"163383e7",
X"f7348452",
X"83e7f451",
X"fe933f83",
X"e0800881",
X"ff068417",
X"33555372",
X"742e8738",
X"fdce3ffe",
X"d13980e4",
X"51ecf13f",
X"873d0d04",
X"f43d0d7e",
X"60595580",
X"5d807582",
X"2b7183ea",
X"94120c83",
X"eaac175b",
X"5b577679",
X"3477772e",
X"83b73876",
X"527751ff",
X"aa943f8e",
X"3dfc0554",
X"905383e9",
X"fc527751",
X"ffa9cf3f",
X"7c567590",
X"2e098106",
X"83933883",
X"e9fc51fc",
X"de3f83e9",
X"fe51fcd7",
X"3f83ea80",
X"51fcd03f",
X"7683ea8c",
X"0c7751ff",
X"a79b3f80",
X"f8885283",
X"e0800851",
X"c9b53f83",
X"e0800881",
X"2e098106",
X"80d43876",
X"83eaa40c",
X"820b83e9",
X"fc34ff96",
X"0b83e9fd",
X"347751ff",
X"a9e13f83",
X"e0800855",
X"83e08008",
X"77258838",
X"83e08008",
X"8f055574",
X"842c7083",
X"ffff0670",
X"882a5851",
X"557583e9",
X"fe347483",
X"e9ff3476",
X"83ea8034",
X"ff800b83",
X"ea813481",
X"903983e9",
X"fc3383e9",
X"fd337188",
X"2b07565b",
X"7483ffff",
X"2e098106",
X"80e838fe",
X"800b83ea",
X"a40c810b",
X"83ea8c0c",
X"ff0b83e9",
X"fc34ff0b",
X"83e9fd34",
X"7751ffa8",
X"ee3f83e0",
X"800883ea",
X"b00c83e0",
X"80085583",
X"e0800880",
X"25883883",
X"e080088f",
X"05557484",
X"2c7083ff",
X"ff067088",
X"2a585155",
X"7583e9fe",
X"347483e9",
X"ff347683",
X"ea8034ff",
X"800b83ea",
X"8134810b",
X"83ea8b34",
X"a5397485",
X"962e0981",
X"0680fe38",
X"7583eaa4",
X"0c7751ff",
X"a8a23f83",
X"ea8b3383",
X"e0800807",
X"557483ea",
X"8b3483ea",
X"8b338106",
X"5574802e",
X"83388457",
X"83ea8033",
X"83ea8133",
X"71882b07",
X"565c7481",
X"802e0981",
X"06a13883",
X"e9fe3383",
X"e9ff3371",
X"882b0756",
X"5bad8075",
X"27873876",
X"8207579c",
X"39768107",
X"57963974",
X"82802e09",
X"81068738",
X"76830757",
X"87397481",
X"ff268a38",
X"7783ea94",
X"1b0c7679",
X"348e3d0d",
X"04803d0d",
X"72842983",
X"ea940570",
X"0883e080",
X"0c51823d",
X"0d04803d",
X"0d727083",
X"e7ec0c70",
X"842980fd",
X"ec057008",
X"83eaa80c",
X"5151823d",
X"0d04fe3d",
X"0d8151de",
X"3f800b83",
X"e9f80c80",
X"0b83e9f4",
X"0cff0b83",
X"e7f00ca8",
X"0b83ea90",
X"0cae51cd",
X"ba3f800b",
X"83ea9454",
X"52807370",
X"8405550c",
X"81125271",
X"842e0981",
X"06ef3884",
X"3d0d04fe",
X"3d0d7402",
X"84059605",
X"22535371",
X"802e9638",
X"72708105",
X"543351cd",
X"c53fff12",
X"7083ffff",
X"065152e7",
X"39843d0d",
X"04fe3d0d",
X"02920522",
X"5382ac51",
X"e7e63f80",
X"c351cda2",
X"3f819651",
X"e7da3f72",
X"5283e7f4",
X"51ffb43f",
X"725283e7",
X"f451f8cd",
X"3f83e080",
X"0881ff06",
X"51ccff3f",
X"843d0d04",
X"ffb13d0d",
X"80d13df8",
X"0551f8f7",
X"3f83e9f8",
X"08810583",
X"e9f80c80",
X"cf3d33cf",
X"117081ff",
X"06515656",
X"74832688",
X"e638758f",
X"06ff0556",
X"7583e7f0",
X"082e9b38",
X"75832696",
X"387583e7",
X"f00c7584",
X"2983ea94",
X"05700853",
X"557551f9",
X"fb3f8076",
X"2488c238",
X"75842983",
X"ea940555",
X"7408802e",
X"88b33883",
X"e7f00884",
X"2983ea94",
X"05700802",
X"880582b9",
X"0533525b",
X"557480d2",
X"2e84b038",
X"7480d224",
X"903874bf",
X"2e9c3874",
X"80d02e81",
X"d53887f2",
X"397480d3",
X"2e80d338",
X"7480d72e",
X"81c43887",
X"e1390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"56cbfb3f",
X"80c151cb",
X"b53ff698",
X"3f83eaab",
X"3383e7f4",
X"34815283",
X"e7f451cc",
X"d23f8151",
X"fde73f74",
X"8b3883ea",
X"a80883ea",
X"900c8739",
X"a80b83ea",
X"900ccbc6",
X"3f80c151",
X"cb803ff5",
X"e33f900b",
X"83ea8b33",
X"81065656",
X"74802e83",
X"38985683",
X"ea803383",
X"ea813371",
X"882b0756",
X"59748180",
X"2e098106",
X"9c3883e9",
X"fe3383e9",
X"ff337188",
X"2b075657",
X"ad807527",
X"8c387581",
X"80075685",
X"3975a007",
X"567583e7",
X"f434ff0b",
X"83e7f534",
X"e00b83e7",
X"f634800b",
X"83e7f734",
X"845283e7",
X"f451cbc7",
X"3f845186",
X"9b390282",
X"bb053302",
X"840582ba",
X"05337182",
X"80290556",
X"59cabb3f",
X"7951ffa2",
X"cf3f83e0",
X"8008802e",
X"8a3880ce",
X"51c9e73f",
X"85f13980",
X"c151c9de",
X"3fcacf3f",
X"c9883f83",
X"eaa40858",
X"8375259b",
X"3883ea80",
X"3383ea81",
X"3371882b",
X"07fc1771",
X"297a0583",
X"80055a51",
X"578d3974",
X"81802918",
X"ff800558",
X"81805780",
X"5676762e",
X"9238c9ba",
X"3f83e080",
X"0883e7f4",
X"17348116",
X"56eb39c9",
X"a93f83e0",
X"800881ff",
X"06775383",
X"e7f45256",
X"f4bf3f83",
X"e0800881",
X"ff065575",
X"752e0981",
X"06819538",
X"9451e3a4",
X"3fc9a33f",
X"80c151c8",
X"dd3fc9ce",
X"3f775279",
X"51ffa0e2",
X"3f805e80",
X"d13dfdf4",
X"05547653",
X"83e7f452",
X"7951ff9e",
X"ef3f0282",
X"b9053355",
X"81597480",
X"d72e0981",
X"0680c538",
X"77527951",
X"ffa0b33f",
X"80d13dfd",
X"f0055476",
X"538f3d70",
X"537a5258",
X"ff9feb3f",
X"80567676",
X"2ea23875",
X"1883e7f4",
X"17337133",
X"70723270",
X"30708025",
X"70307f06",
X"811d5d5f",
X"51515152",
X"5b55db39",
X"82ac51e2",
X"9f3f7880",
X"2e863880",
X"c3518439",
X"80ce51c7",
X"d13fc8c2",
X"3fc6fb3f",
X"83d83902",
X"82bb0533",
X"02840582",
X"ba053371",
X"82802905",
X"59558070",
X"5d5980e4",
X"51e1e93f",
X"c7e83f80",
X"c151c7a2",
X"3f83ea8c",
X"08792e82",
X"d63883ea",
X"b00880fc",
X"055580fd",
X"52745185",
X"c13f83e0",
X"80085b77",
X"8224b238",
X"ff187087",
X"2b83ffff",
X"800680fc",
X"b80583e7",
X"f4595755",
X"81805575",
X"70810557",
X"33777081",
X"055934ff",
X"157081ff",
X"06515574",
X"ea388285",
X"397782e8",
X"2e81a338",
X"7782e92e",
X"09810681",
X"aa387858",
X"77873270",
X"30707207",
X"80257a8a",
X"32703070",
X"72078025",
X"73075354",
X"5a515755",
X"75802e97",
X"38787826",
X"9238a00b",
X"83e7f41a",
X"34811970",
X"81ff065a",
X"55eb3981",
X"187081ff",
X"0659558a",
X"7827ffbc",
X"388f5883",
X"e7ef1833",
X"83e7f419",
X"34ff1870",
X"81ff0659",
X"55778426",
X"ea389058",
X"800b83e7",
X"f4193481",
X"187081ff",
X"0670982b",
X"52595574",
X"8025e938",
X"80c6557a",
X"858f2484",
X"3880c255",
X"7483e7f4",
X"3480f10b",
X"83e7f734",
X"810b83e7",
X"f8347a83",
X"e7f5347a",
X"882c5574",
X"83e7f634",
X"80cb3982",
X"f0782580",
X"c4387780",
X"fd29fd97",
X"d3055279",
X"51ff9d8e",
X"3f80d13d",
X"fdec0554",
X"80fd5383",
X"e7f45279",
X"51ff9cc6",
X"3f7b8119",
X"59567580",
X"fc248338",
X"78587788",
X"2c557483",
X"e8f13477",
X"83e8f234",
X"7583e8f3",
X"34818059",
X"80cc3983",
X"eaa40857",
X"8378259b",
X"3883ea80",
X"3383ea81",
X"3371882b",
X"07fc1a71",
X"29790583",
X"80055951",
X"598d3977",
X"81802917",
X"ff800557",
X"81805976",
X"527951ff",
X"9c9c3f80",
X"d13dfdec",
X"05547853",
X"83e7f452",
X"7951ff9b",
X"d53f7851",
X"f6bf3fc4",
X"e53fc39e",
X"3f8b3983",
X"e9f40881",
X"0583e9f4",
X"0c80d13d",
X"0d04f6e0",
X"3ffc39fc",
X"3d0d7678",
X"71842983",
X"ea940570",
X"08515353",
X"53709e38",
X"80ce7234",
X"80cf0b81",
X"133480ce",
X"0b821334",
X"80c50b83",
X"13347084",
X"133480e7",
X"3983eaac",
X"13335480",
X"d2723473",
X"822a7081",
X"06515180",
X"cf537084",
X"3880d753",
X"72811334",
X"a00b8213",
X"34738306",
X"5170812e",
X"9e387081",
X"24883870",
X"802e8f38",
X"9f397082",
X"2e923870",
X"832e9238",
X"933980d8",
X"558e3980",
X"d3558939",
X"80cd5584",
X"3980c455",
X"74831334",
X"80c40b84",
X"1334800b",
X"85133486",
X"3d0d0483",
X"e7ec0883",
X"e0800c04",
X"803d0d83",
X"e7ec0884",
X"2980fe8c",
X"05700883",
X"e0800c51",
X"823d0d04",
X"fc3d0d76",
X"78535481",
X"53805587",
X"39711073",
X"10545273",
X"72265172",
X"802ea738",
X"70802e86",
X"38718025",
X"e8387280",
X"2e983871",
X"74268938",
X"73723175",
X"74075654",
X"72812a72",
X"812a5353",
X"e5397351",
X"78833874",
X"517083e0",
X"800c863d",
X"0d04fe3d",
X"0d805375",
X"527451ff",
X"a33f843d",
X"0d04fe3d",
X"0d815375",
X"527451ff",
X"933f843d",
X"0d04fb3d",
X"0d777955",
X"55805674",
X"76258638",
X"74305581",
X"56738025",
X"88387330",
X"76813257",
X"54805373",
X"527451fe",
X"e73f83e0",
X"80085475",
X"802e8738",
X"83e08008",
X"30547383",
X"e0800c87",
X"3d0d04fa",
X"3d0d787a",
X"57558057",
X"74772586",
X"38743055",
X"8157759f",
X"2c548153",
X"75743274",
X"31527451",
X"feaa3f83",
X"e0800854",
X"76802e87",
X"3883e080",
X"08305473",
X"83e0800c",
X"883d0d04",
X"fd3d0d75",
X"5480740c",
X"800b8415",
X"0c800b88",
X"150c800b",
X"8c150c87",
X"a6803370",
X"81ff0670",
X"71842a06",
X"515151da",
X"aa3f7081",
X"2a813271",
X"81327181",
X"06718106",
X"3184170c",
X"53537083",
X"2a813271",
X"822a8132",
X"70810672",
X"7131770c",
X"51525287",
X"a0903387",
X"a0913370",
X"81ff0670",
X"73068132",
X"81068818",
X"0c515252",
X"83e08008",
X"802e80c2",
X"3883e080",
X"08812a70",
X"810683e0",
X"80088106",
X"3184160c",
X"5183e080",
X"08832a83",
X"e0800882",
X"2a718106",
X"71810631",
X"760c5252",
X"83e08008",
X"842a8106",
X"88150c83",
X"e0800885",
X"2a81068c",
X"150c853d",
X"0d04fe3d",
X"0d747654",
X"527151fe",
X"bb3f7281",
X"2ea23881",
X"73268d38",
X"72822ea8",
X"3872832e",
X"9c38e639",
X"7108e238",
X"841208dd",
X"38881208",
X"d838a539",
X"88120881",
X"2e9e3891",
X"39881208",
X"812e9538",
X"71089138",
X"8412088c",
X"388c1208",
X"812e0981",
X"06ffb238",
X"843d0d04",
X"00ffffff",
X"ff00ffff",
X"ffff00ff",
X"ffffff00",
X"809a9041",
X"8e418f80",
X"45454549",
X"49498e8f",
X"9092924f",
X"994f5555",
X"59999a9b",
X"9c9d9e9f",
X"41494f55",
X"a5a5a6a7",
X"a8a9aaab",
X"ac21aeaf",
X"b0b1b2b3",
X"b4b5b6b7",
X"b8b9babb",
X"bcbdbebf",
X"c0c1c2c3",
X"c4c5c6c7",
X"c8c9cacb",
X"cccdcecf",
X"d0d1d2d3",
X"d4d5d6d7",
X"d8d9dadb",
X"dcdddedf",
X"e0e1e2e3",
X"e4e5e6e7",
X"e8e9eaeb",
X"ecedeeef",
X"f0f1f2f3",
X"f4f5f6f7",
X"f8f9fafb",
X"fcfdfeff",
X"00002bd4",
X"00002c15",
X"00002c37",
X"00002c59",
X"00002c7f",
X"00002c7f",
X"00002c7f",
X"00002c7f",
X"00002cf0",
X"00002d45",
X"00002d45",
X"00002d85",
X"2e2e0000",
X"25732025",
X"73000000",
X"20000000",
X"41545200",
X"58464400",
X"58455800",
X"43686f6f",
X"73652000",
X"66696c65",
X"00000000",
X"4449523a",
X"00000000",
X"44495200",
X"25303278",
X"00000000",
X"36344b00",
X"3132384b",
X"00000000",
X"3332304b",
X"28436f6d",
X"70792900",
X"3332304b",
X"2852616d",
X"626f2900",
X"3537364b",
X"28436f6d",
X"70792900",
X"3537364b",
X"2852616d",
X"626f2900",
X"314d4200",
X"344d4200",
X"53650000",
X"7474696e",
X"67730000",
X"43505520",
X"54757262",
X"6f3a2564",
X"78000000",
X"44726976",
X"65205475",
X"72626f3a",
X"25730000",
X"52616d3a",
X"25730000",
X"526f6d3a",
X"25730000",
X"44726976",
X"65202564",
X"3a257320",
X"25730000",
X"4e4f4e45",
X"00000000",
X"43617274",
X"3a202573",
X"00000000",
X"4c6f6164",
X"206d656d",
X"6f727900",
X"53617665",
X"206d656d",
X"6f727920",
X"28666f72",
X"20646562",
X"75676769",
X"6e672900",
X"45786974",
X"00000000",
X"61746172",
X"69626173",
X"2e726f6d",
X"00000000",
X"61746172",
X"69786c2e",
X"726f6d00",
X"524f4d00",
X"42494e00",
X"43415200",
X"4d454d00",
X"5374616e",
X"64617264",
X"00000000",
X"46617374",
X"28362900",
X"46617374",
X"28352900",
X"46617374",
X"28342900",
X"46617374",
X"28332900",
X"46617374",
X"28322900",
X"46617374",
X"28312900",
X"46617374",
X"28302900",
X"00000000",
X"00000000",
X"01010008",
X"02210010",
X"080d0040",
X"090a0040",
X"0a090040",
X"0b080040",
X"0c300020",
X"0d310040",
X"0e320080",
X"0f040010",
X"110c0080",
X"17330100",
X"18340200",
X"1a280010",
X"1b290020",
X"1c2a0040",
X"1d2b0080",
X"1e2c0100",
X"1f2d0200",
X"21380020",
X"22390040",
X"233a0080",
X"243b0100",
X"253c0200",
X"28230010",
X"29020080",
X"2a030400",
X"38240200",
X"00000000",
X"70704740",
X"2c704268",
X"2c020202",
X"02020202",
X"02020202",
X"02020202",
X"02020202",
X"02020241",
X"00060000",
X"00003c34",
X"00003c38",
X"00003c40",
X"00003c4c",
X"00003c58",
X"00003c64",
X"00003c70",
X"00003c74",
X"72025f07",
X"f807a900",
X"8d04038d",
X"4402a907",
X"8d0503a9",
X"708d0a03",
X"a9018d0b",
X"03850960",
X"7d8a4820",
X"53e488d0",
X"fa68aa8c",
X"8e07ad7d",
X"07ee8e07",
X"60a9938d",
X"e202a907",
X"8de302a2",
X"0220da07",
X"954320da",
X"07954435",
X"43c9fff0",
X"f0caca10",
X"ec3006e6",
X"45d002e6",
X"4620da07",
X"a2018144",
X"b545d543",
X"d0edca10",
X"f720d207",
X"4c9407a9",
X"038d0fd2",
X"6ce202ad",
X"8e07cd7f",
X"07d0abee",
X"0a03d003",
X"ee0b03ad",
X"7d070d7e",
X"07d08e20",
X"d2076ce0",
X"0220da07",
X"8de00220",
X"da078de1",
X"022de002",
X"c9fff0ed",
X"a9008d8e",
X"07f08200",
X"00000028",
X"00000006",
X"00000005",
X"00000004",
X"00000003",
X"00000002",
X"00000001",
X"00000000",
X"00003d34",
X"00003d40",
X"00003d48",
X"00003d50",
X"00003d58",
X"00003d60",
X"00003d68",
X"00003d70",
X"2f617461",
X"72693830",
X"302f726f",
X"6d000000",
X"2f617461",
X"72693830",
X"302f7573",
X"65720000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000",
X"00000000"

);
        signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
