-------------------------------------------------------------------------------
--
-- SNESpad controller core
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- $Id: snespad_pad-c.vhd,v 1.1 2004/10/05 17:01:27 arniml Exp $
--
-------------------------------------------------------------------------------

configuration snespad_pad_rtl_c0 of snespad_pad is

  for rtl
  end for;

end snespad_pad_rtl_c0;
