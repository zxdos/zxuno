library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity PointerRamBlack is

    port (
        clka  : in  std_logic;
        wea   : in  std_logic;
        addra : in  std_logic_vector(7 downto 0);
        dina  : in  std_logic_vector(7 downto 0);
        douta : out std_logic_vector(7 downto 0);
        clkb  : in  std_logic;
        web   : in  std_logic;
        addrb : in  std_logic_vector(7 downto 0);
        dinb  : in  std_logic_vector(7 downto 0);
        doutb : out std_logic_vector(7 downto 0)
        );
end PointerRamBlack;

architecture BEHAVIORAL of PointerRamBlack is

-- Shared memory
    type ram_type is array (0 to 255) of std_logic_vector (7 downto 0);
    shared variable RAM : ram_type := (
        "11111111",
        "10000010",
        "10000100",
        "10000100",
        "10000010",
        "10110001",
        "11001010",
        "10000100",

        "11100000",
        "10100000",
        "11100000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",

        "00111100",
        "01010010",
        "10010001",
        "10010001",
        "10011101",
        "10000001",
        "01000010",
        "00111100",

        "11111111",
        "10000001",
        "10111111",
        "10100000",
        "10100000",
        "10100000",
        "10100000",
        "11100000",

        "00010000",
        "00101000",
        "01000100",
        "11000110",
        "01000100",
        "01000100",
        "01000100",
        "01111100",

        "01111100",
        "01000100",
        "01000100",
        "01000100",
        "11000110",
        "01000100",
        "00101000",
        "00010000",

        "00001000",
        "11111100",
        "10000010",
        "10000001",
        "10000010",
        "11111100",
        "00001000",
        "00000000",

        "00010000",
        "00111111",
        "01000001",
        "10000001",
        "01000001",
        "00111111",
        "00010000",
        "00000000",

        "00111100",
        "01000110",
        "10001101",
        "10001101",
        "10011001",
        "10011001",
        "01110010",
        "00111100",

        "00111000",
        "01000100",
        "01010100",
        "01110100",
        "00101000",
        "00111000",
        "00101000",
        "00111000",

        "01111100",
        "01000100",
        "01101100",
        "00101000",
        "00101000",
        "01101100",
        "01000100",
        "01111100",

        "00111000",
        "00101000",
        "11101110",
        "10000010",
        "11101110",
        "00101000",
        "00111000",
        "00000000",

        "01000000",
        "10100000",
        "10100000",
        "10111110",
        "10101011",
        "10000001",
        "11111111",
        "01111110",

        "01111110",
        "11111111",
        "10000001",
        "10101011",
        "10111110",
        "10100000",
        "10100000",
        "01000000",

        "01111110",
        "11000001",
        "11011110",
        "11001000",
        "11011000",
        "11001000",
        "11011000",
        "01110000",

        "01111110",
        "10000011",
        "01111011",
        "00010011",
        "00011011",
        "00010011",
        "00011011",
        "00001110",

        "11111111",
        "01000010",
        "00100100",
        "00011000",
        "00011000",
        "00100100",
        "01000010",
        "11111111",

        "11111111",
        "01000010",
        "00100100",
        "00011000",
        "00011000",
        "00100100",
        "01011010",
        "11111111",

        "11111111",
        "01000010",
        "00100100",
        "00011000",
        "00011000",
        "00100100",
        "01111110",
        "11111111",

        "11111111",
        "01000010",
        "00100100",
        "00011000",
        "00011000",
        "00111100",
        "01111110",
        "11111111",

        "11100000",
        "10011000",
        "01000110",
        "00110001",
        "01101011",
        "01010101",
        "00101001",
        "00011110",

        "00000111",
        "00011001",
        "01100010",
        "10001100",
        "11010110",
        "10101010",
        "10010100",
        "01111000",

        "00011110",
        "00101001",
        "01010101",
        "01101011",
        "00110001",
        "01000110",
        "10011000",
        "11100000",

        "01111000",
        "10010100",
        "10101010",
        "11010110",
        "10001100",
        "01100010",
        "00011001",
        "00000111",

        "01100110",
        "10011001",
        "10011001",
        "11011101",
        "11011101",
        "10011001",
        "10011001",
        "01100110",

        "01100110",
        "11111111",
        "11111111",
        "10011001",
        "10011001",
        "10011001",
        "10011001",
        "01100110",

        "01100110",
        "10011001",
        "10011001",
        "10111011",
        "10111011",
        "10011001",
        "10011001",
        "01100110",

        "01100110",
        "10011001",
        "10011001",
        "10011001",
        "10011001",
        "11111111",
        "11111111",
        "01100110",

        "11111111",
        "10000010",
        "10000100",
        "10001000",
        "10010000",
        "10100000",
        "11000000",
        "10000000",

        "10000000",
        "11000000",
        "10100000",
        "10010000",
        "10001000",
        "10000100",
        "10000010",
        "11111111",

        "00000001",
        "00000011",
        "00000101",
        "00001001",
        "00010001",
        "00100001",
        "01000001",
        "11111111",

        "11111111",
        "01000001",
        "00100001",
        "00010001",
        "00001001",
        "00000101",
        "00000011",
        "00000001"
        );

--attribute RAM_STYLE : string;
--attribute RAM_STYLE of RAM: signal is "BLOCK";

begin

    process (clka)
    begin
        if rising_edge(clka) then
            if (wea = '1') then
                RAM(conv_integer(addra(7 downto 0))) := dina;
            end if;
            douta <= RAM(conv_integer(addra(7 downto 0)));
        end if;
    end process;

    process (clkb)
    begin
        if rising_edge(clkb) then
            if (web = '1') then
                RAM(conv_integer(addrb(7 downto 0))) := dinb;
            end if;
            doutb <= RAM(conv_integer(addrb(7 downto 0)));
        end if;
    end process;

end BEHAVIORAL;

