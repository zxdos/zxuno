
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity os16_loop is
port(
        clock:in std_logic;
        address:in std_logic_vector(13 downto 0);
        q:out std_logic_vector(7 downto 0)
);
end os16_loop;

architecture syn of os16_loop is
        type rom_type is array(0 to 16383) of std_logic_vector(7 downto 0);
        signal ROM:rom_type:=
(
X"a9", --X"a2", -- LDX
X"12", --X"00",
X"8d", --X"e8",
X"01", --X"8a",
X"00", --X"8d",
X"a9", --X"10",
X"34", --X"00",
X"8d", --X"ad",
--
X"02", --X"10",
X"00", --X"00",
X"a9", --X"4c",
X"56", --X"02",
X"8d", --X"c0",
X"03", --X"40",
X"00", --X"8d",
X"a9", --X"0e",
--
X"67", --X"d4",
X"8d", --X"ad",
X"04", --X"13",
X"00", --X"d0",
X"ad", --X"8d",
X"01", --X"fa",
X"00", --X"03",
X"ad", --X"60",
--
X"02", --X"2c",
X"00", --X"0f",
X"ad", --X"d4",
X"03", --X"10",
X"00", --X"03",
X"ad", --X"6c",
X"04", --X"00",
X"00", --X"02",

X"4c", --X"d8",
X"00", --X"48",
X"c0", --X"8a",

X"48",
X"98",
X"48",
X"8d",
X"0f",
X"d4",
X"6c",
X"22",
X"02",
X"d8",
X"6c",
X"16",
X"02",
X"48",
X"ad",
X"0e",
X"d2",
X"29",
X"20",
X"d0",
X"0d",
X"a9",
X"df",
X"8d",
X"0e",
X"d2",
X"a5",
X"10",
X"8d",
X"0e",
X"d2",
X"6c",
X"0a",
X"02",
X"8a",
X"48",
X"ad",
X"ff",
X"d1",
X"2d",
X"49",
X"02",
X"f0",
X"03",
X"6c",
X"38",
X"02",
X"a2",
X"06",
X"bd",
X"cf",
X"c0",
X"e0",
X"05",
X"d0",
X"04",
X"25",
X"10",
X"f0",
X"05",
X"2c",
X"0e",
X"d2",
X"f0",
X"06",
X"ca",
X"10",
X"ed",
X"4c",
X"a0",
X"c0",
X"49",
X"ff",
X"8d",
X"0e",
X"d2",
X"a5",
X"10",
X"8d",
X"0e",
X"d2",
X"e0",
X"00",
X"d0",
X"05",
X"ad",
X"6d",
X"02",
X"d0",
X"23",
X"bd",
X"d7",
X"c0",
X"aa",
X"bd",
X"00",
X"02",
X"8d",
X"8c",
X"02",
X"bd",
X"01",
X"02",
X"8d",
X"8d",
X"02",
X"68",
X"aa",
X"6c",
X"8c",
X"02",
X"a9",
X"00",
X"85",
X"11",
X"8d",
X"ff",
X"02",
X"8d",
X"f0",
X"02",
X"85",
X"4d",
X"68",
X"40",
X"68",
X"aa",
X"2c",
X"02",
X"d3",
X"10",
X"06",
X"ad",
X"00",
X"d3",
X"6c",
X"02",
X"02",
X"2c",
X"03",
X"d3",
X"10",
X"06",
X"ad",
X"01",
X"d3",
X"6c",
X"04",
X"02",
X"68",
X"8d",
X"8c",
X"02",
X"68",
X"48",
X"29",
X"10",
X"f0",
X"07",
X"ad",
X"8c",
X"02",
X"48",
X"6c",
X"06",
X"02",
X"ad",
X"8c",
X"02",
X"48",
X"68",
X"40",
X"80",
X"40",
X"04",
X"02",
X"01",
X"08",
X"10",
X"20",
X"36",
X"08",
X"14",
X"12",
X"10",
X"0e",
X"0c",
X"0a",
X"4c",
X"df",
X"c0",
X"e6",
X"14",
X"d0",
X"08",
X"e6",
X"4d",
X"e6",
X"13",
X"d0",
X"02",
X"e6",
X"12",
X"a9",
X"fe",
X"a2",
X"00",
X"a4",
X"4d",
X"10",
X"06",
X"85",
X"4d",
X"a6",
X"13",
X"a9",
X"f6",
X"85",
X"4e",
X"86",
X"4f",
X"ad",
X"c5",
X"02",
X"45",
X"4f",
X"25",
X"4e",
X"8d",
X"17",
X"d0",
X"a2",
X"00",
X"20",
X"55",
X"c2",
X"d0",
X"03",
X"20",
X"4f",
X"c2",
X"a5",
X"42",
X"d0",
X"08",
X"ba",
X"bd",
X"04",
X"01",
X"29",
X"04",
X"f0",
X"03",
X"4c",
X"8a",
X"c2",
X"ad",
X"13",
X"d0",
X"cd",
X"fa",
X"03",
X"d0",
X"b4",
X"ad",
X"0d",
X"d4",
X"8d",
X"35",
X"02",
X"ad",
X"0c",
X"d4",
X"8d",
X"34",
X"02",
X"ad",
X"31",
X"02",
X"8d",
X"03",
X"d4",
X"ad",
X"30",
X"02",
X"8d",
X"02",
X"d4",
X"ad",
X"2f",
X"02",
X"8d",
X"00",
X"d4",
X"ad",
X"6f",
X"02",
X"8d",
X"1b",
X"d0",
X"ad",
X"6c",
X"02",
X"f0",
X"0e",
X"ce",
X"6c",
X"02",
X"a9",
X"08",
X"38",
X"ed",
X"6c",
X"02",
X"29",
X"07",
X"8d",
X"05",
X"d4",
X"a2",
X"08",
X"8e",
X"1f",
X"d0",
X"58",
X"bd",
X"c0",
X"02",
X"45",
X"4f",
X"25",
X"4e",
X"9d",
X"12",
X"d0",
X"ca",
X"10",
X"f2",
X"ad",
X"f4",
X"02",
X"8d",
X"09",
X"d4",
X"ad",
X"f3",
X"02",
X"8d",
X"01",
X"d4",
X"a2",
X"02",
X"20",
X"55",
X"c2",
X"d0",
X"03",
X"20",
X"52",
X"c2",
X"a2",
X"02",
X"e8",
X"e8",
X"bd",
X"18",
X"02",
X"1d",
X"19",
X"02",
X"f0",
X"06",
X"20",
X"55",
X"c2",
X"9d",
X"26",
X"02",
X"e0",
X"08",
X"d0",
X"ec",
X"ad",
X"0f",
X"d2",
X"29",
X"04",
X"f0",
X"08",
X"ad",
X"f1",
X"02",
X"f0",
X"03",
X"ce",
X"f1",
X"02",
X"ad",
X"2b",
X"02",
X"f0",
X"3e",
X"ad",
X"0f",
X"d2",
X"29",
X"04",
X"d0",
X"32",
X"ce",
X"2b",
X"02",
X"d0",
X"32",
X"ad",
X"6d",
X"02",
X"d0",
X"2d",
X"ad",
X"da",
X"02",
X"8d",
X"2b",
X"02",
X"ad",
X"09",
X"d2",
X"c9",
X"9f",
X"f0",
X"20",
X"c9",
X"83",
X"f0",
X"1c",
X"c9",
X"84",
X"f0",
X"18",
X"c9",
X"94",
X"f0",
X"14",
X"29",
X"3f",
X"c9",
X"11",
X"f0",
X"0e",
X"ad",
X"09",
X"d2",
X"8d",
X"fc",
X"02",
X"4c",
X"f3",
X"c1",
X"a9",
X"00",
X"8d",
X"2b",
X"02",
X"ad",
X"00",
X"d3",
X"4a",
X"4a",
X"4a",
X"4a",
X"8d",
X"79",
X"02",
X"8d",
X"7b",
X"02",
X"ad",
X"00",
X"d3",
X"29",
X"0f",
X"8d",
X"78",
X"02",
X"8d",
X"7a",
X"02",
X"ad",
X"10",
X"d0",
X"8d",
X"84",
X"02",
X"8d",
X"86",
X"02",
X"ad",
X"11",
X"d0",
X"8d",
X"85",
X"02",
X"8d",
X"87",
X"02",
X"a2",
X"03",
X"bd",
X"00",
X"d2",
X"9d",
X"70",
X"02",
X"9d",
X"74",
X"02",
X"ca",
X"10",
X"f4",
X"8d",
X"0b",
X"d2",
X"a2",
X"02",
X"a0",
X"01",
X"b9",
X"78",
X"02",
X"4a",
X"4a",
X"4a",
X"9d",
X"7d",
X"02",
X"9d",
X"81",
X"02",
X"a9",
X"00",
X"2a",
X"9d",
X"7c",
X"02",
X"9d",
X"80",
X"02",
X"ca",
X"ca",
X"88",
X"10",
X"e6",
X"6c",
X"24",
X"02",
X"6c",
X"26",
X"02",
X"6c",
X"28",
X"02",
X"bc",
X"18",
X"02",
X"d0",
X"08",
X"bc",
X"19",
X"02",
X"f0",
X"10",
X"de",
X"19",
X"02",
X"de",
X"18",
X"02",
X"d0",
X"08",
X"bc",
X"19",
X"02",
X"d0",
X"03",
X"a9",
X"00",
X"60",
X"a9",
X"ff",
X"60",
X"0a",
X"8d",
X"2d",
X"02",
X"8a",
X"a2",
X"05",
X"8d",
X"0a",
X"d4",
X"ca",
X"d0",
X"fd",
X"ae",
X"2d",
X"02",
X"9d",
X"17",
X"02",
X"98",
X"9d",
X"16",
X"02",
X"60",
X"68",
X"a8",
X"68",
X"aa",
X"68",
X"40",
X"78",
X"ad",
X"13",
X"d0",
X"cd",
X"fa",
X"03",
X"d0",
X"2f",
X"6a",
X"90",
X"05",
X"20",
X"c9",
X"c4",
X"d0",
X"27",
X"ad",
X"44",
X"02",
X"d0",
X"22",
X"a9",
X"ff",
X"d0",
X"20",
X"78",
X"a2",
X"8c",
X"88",
X"d0",
X"fd",
X"ca",
X"d0",
X"fa",
X"ad",
X"3d",
X"03",
X"c9",
X"5c",
X"d0",
X"0e",
X"ad",
X"3e",
X"03",
X"c9",
X"93",
X"d0",
X"07",
X"ad",
X"3f",
X"03",
X"c9",
X"25",
X"f0",
X"c8",
X"a9",
X"00",
X"85",
X"08",
X"78",
X"d8",
X"a2",
X"ff",
X"9a",
X"20",
X"71",
X"c4",
X"a9",
X"01",
X"85",
X"01",
X"a5",
X"08",
X"d0",
X"52",
X"a9",
X"00",
X"a0",
X"08",
X"85",
X"04",
X"85",
X"05",
X"a9",
X"ff",
X"91",
X"04",
X"d1",
X"04",
X"f0",
X"02",
X"46",
X"01",
X"a9",
X"00",
X"91",
X"04",
X"d1",
X"04",
X"f0",
X"02",
X"46",
X"01",
X"c8",
X"d0",
X"e9",
X"e6",
X"05",
X"a6",
X"05",
X"e4",
X"06",
X"d0",
X"e1",
X"a9",
X"23",
X"85",
X"0a",
X"a9",
X"f2",
X"85",
X"0b",
X"ad",
X"01",
X"d3",
X"29",
X"7f",
X"8d",
X"01",
X"d3",
X"20",
X"73",
X"ff",
X"b0",
X"05",
X"20",
X"92",
X"ff",
X"90",
X"02",
X"46",
X"01",
X"ad",
X"01",
X"d3",
X"09",
X"80",
X"8d",
X"01",
X"d3",
X"a9",
X"ff",
X"8d",
X"44",
X"02",
X"d0",
X"22",
X"a2",
X"00",
X"ad",
X"ec",
X"03",
X"f0",
X"07",
X"8e",
X"0e",
X"00",
X"8e",
X"0f",
X"00",
X"8a",
X"9d",
X"00",
X"02",
X"e0",
X"ed",
X"b0",
X"03",
X"9d",
X"00",
X"03",
X"ca",
X"d0",
X"f3",
X"a2",
X"10",
X"95",
X"00",
X"e8",
X"10",
X"fb",
X"a2",
X"00",
X"ad",
X"01",
X"d3",
X"29",
X"02",
X"f0",
X"01",
X"e8",
X"8e",
X"f8",
X"03",
X"a9",
X"5c",
X"8d",
X"3d",
X"03",
X"a9",
X"93",
X"8d",
X"3e",
X"03",
X"a9",
X"25",
X"8d",
X"3f",
X"03",
X"a9",
X"02",
X"85",
X"52",
X"a9",
X"27",
X"85",
X"53",
X"ad",
X"14",
X"d0",
X"29",
X"0e",
X"d0",
X"08",
X"a9",
X"05",
X"a2",
X"01",
X"a0",
X"28",
X"d0",
X"06",
X"a9",
X"06",
X"a2",
X"00",
X"a0",
X"30",
X"8d",
X"da",
X"02",
X"86",
X"62",
X"8c",
X"d9",
X"02",
X"a2",
X"25",
X"bd",
X"4b",
X"c4",
X"9d",
X"00",
X"02",
X"ca",
X"10",
X"f7",
X"a2",
X"0e",
X"bd",
X"2e",
X"c4",
X"9d",
X"1a",
X"03",
X"ca",
X"10",
X"f7",
X"20",
X"35",
X"c5",
X"58",
X"a5",
X"01",
X"d0",
X"15",
X"ad",
X"01",
X"d3",
X"29",
X"7f",
X"8d",
X"01",
X"d3",
X"a9",
X"02",
X"8d",
X"f3",
X"02",
X"a9",
X"e0",
X"8d",
X"f4",
X"02",
X"4c",
X"03",
X"50",
X"a2",
X"00",
X"86",
X"06",
X"ae",
X"e4",
X"02",
X"e0",
X"b0",
X"b0",
X"0d",
X"ae",
X"fc",
X"bf",
X"d0",
X"08",
X"e6",
X"06",
X"20",
X"c9",
X"c4",
X"20",
X"29",
X"c4",
X"a9",
X"03",
X"a2",
X"00",
X"9d",
X"42",
X"03",
X"a9",
X"48",
X"9d",
X"44",
X"03",
X"a9",
X"c4",
X"9d",
X"45",
X"03",
X"a9",
X"0c",
X"9d",
X"4a",
X"03",
X"20",
X"56",
X"e4",
X"10",
X"03",
X"4c",
X"aa",
X"c2",
X"e8",
X"d0",
X"fd",
X"c8",
X"10",
X"fa",
X"20",
X"6e",
X"c6",
X"a5",
X"06",
X"f0",
X"06",
X"ad",
X"fd",
X"bf",
X"6a",
X"90",
X"06",
X"20",
X"8b",
X"c5",
X"20",
X"39",
X"e7",
X"a9",
X"00",
X"8d",
X"44",
X"02",
X"a5",
X"06",
X"f0",
X"0a",
X"ad",
X"fd",
X"bf",
X"29",
X"04",
X"f0",
X"03",
X"6c",
X"fa",
X"bf",
X"6c",
X"0a",
X"00",
X"6c",
X"fe",
X"bf",
X"18",
X"60",
X"50",
X"30",
X"e4",
X"43",
X"40",
X"e4",
X"45",
X"00",
X"e4",
X"53",
X"10",
X"e4",
X"4b",
X"20",
X"e4",
X"42",
X"4f",
X"4f",
X"54",
X"20",
X"45",
X"52",
X"52",
X"4f",
X"52",
X"9b",
X"45",
X"3a",
X"9b",
X"ce",
X"c0",
X"cd",
X"c0",
X"cd",
X"c0",
X"cd",
X"c0",
X"19",
X"fc",
X"2c",
X"eb",
X"ad",
X"ea",
X"ec",
X"ea",
X"cd",
X"c0",
X"cd",
X"c0",
X"cd",
X"c0",
X"30",
X"c0",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"e2",
X"c0",
X"8a",
X"c2",
X"ad",
X"13",
X"d0",
X"6a",
X"90",
X"0d",
X"ad",
X"fc",
X"bf",
X"d0",
X"08",
X"ad",
X"fd",
X"bf",
X"10",
X"03",
X"6c",
X"fe",
X"bf",
X"20",
X"da",
X"c4",
X"ad",
X"01",
X"d3",
X"09",
X"02",
X"8d",
X"01",
X"d3",
X"a5",
X"08",
X"f0",
X"07",
X"ad",
X"f8",
X"03",
X"d0",
X"11",
X"f0",
X"07",
X"ad",
X"1f",
X"d0",
X"29",
X"04",
X"f0",
X"08",
X"ad",
X"01",
X"d3",
X"29",
X"fd",
X"8d",
X"01",
X"d3",
X"a9",
X"00",
X"a8",
X"85",
X"05",
X"a9",
X"28",
X"85",
X"06",
X"b1",
X"05",
X"49",
X"ff",
X"91",
X"05",
X"d1",
X"05",
X"d0",
X"0c",
X"49",
X"ff",
X"91",
X"05",
X"d1",
X"05",
X"d0",
X"04",
X"e6",
X"06",
X"d0",
X"ea",
X"60",
X"a9",
X"00",
X"aa",
X"18",
X"7d",
X"f0",
X"bf",
X"e8",
X"d0",
X"fa",
X"cd",
X"eb",
X"03",
X"8d",
X"eb",
X"03",
X"60",
X"a9",
X"00",
X"aa",
X"8d",
X"03",
X"d3",
X"9d",
X"00",
X"d0",
X"9d",
X"00",
X"d4",
X"9d",
X"00",
X"d2",
X"e0",
X"01",
X"f0",
X"03",
X"9d",
X"00",
X"d3",
X"e8",
X"d0",
X"ed",
X"a9",
X"3c",
X"8d",
X"03",
X"d3",
X"a9",
X"ff",
X"8d",
X"01",
X"d3",
X"a9",
X"38",
X"8d",
X"02",
X"d3",
X"8d",
X"03",
X"d3",
X"a9",
X"00",
X"8d",
X"00",
X"d3",
X"a9",
X"ff",
X"8d",
X"01",
X"d3",
X"a9",
X"3c",
X"8d",
X"02",
X"d3",
X"8d",
X"03",
X"d3",
X"ad",
X"01",
X"d3",
X"ad",
X"00",
X"d3",
X"a9",
X"22",
X"8d",
X"0f",
X"d2",
X"a9",
X"a0",
X"8d",
X"05",
X"d2",
X"8d",
X"07",
X"d2",
X"a9",
X"28",
X"8d",
X"08",
X"d2",
X"a9",
X"ff",
X"8d",
X"0d",
X"d2",
X"60",
X"c6",
X"11",
X"a9",
X"92",
X"8d",
X"36",
X"02",
X"a9",
X"c0",
X"8d",
X"37",
X"02",
X"a5",
X"06",
X"8d",
X"e4",
X"02",
X"8d",
X"e6",
X"02",
X"a9",
X"00",
X"8d",
X"e5",
X"02",
X"a9",
X"00",
X"8d",
X"e7",
X"02",
X"a9",
X"07",
X"8d",
X"e8",
X"02",
X"20",
X"0c",
X"e4",
X"20",
X"1c",
X"e4",
X"20",
X"2c",
X"e4",
X"20",
X"3c",
X"e4",
X"20",
X"4c",
X"e4",
X"20",
X"6e",
X"e4",
X"20",
X"65",
X"e4",
X"20",
X"6b",
X"e4",
X"20",
X"50",
X"e4",
X"a9",
X"6e",
X"8d",
X"38",
X"02",
X"a9",
X"c9",
X"8d",
X"39",
X"02",
X"20",
X"9b",
X"e4",
X"ad",
X"1f",
X"d0",
X"29",
X"01",
X"49",
X"01",
X"8d",
X"e9",
X"03",
X"60",
X"a5",
X"08",
X"f0",
X"09",
X"a5",
X"09",
X"29",
X"01",
X"f0",
X"33",
X"4c",
X"3b",
X"c6",
X"a9",
X"01",
X"8d",
X"01",
X"03",
X"a9",
X"53",
X"8d",
X"02",
X"03",
X"20",
X"53",
X"e4",
X"30",
X"21",
X"a9",
X"00",
X"8d",
X"0b",
X"03",
X"a9",
X"01",
X"8d",
X"0a",
X"03",
X"a9",
X"00",
X"8d",
X"04",
X"03",
X"a9",
X"04",
X"8d",
X"05",
X"03",
X"20",
X"59",
X"c6",
X"10",
X"09",
X"20",
X"3e",
X"c6",
X"ad",
X"ea",
X"03",
X"f0",
X"df",
X"60",
X"a2",
X"03",
X"bd",
X"00",
X"04",
X"9d",
X"40",
X"02",
X"ca",
X"10",
X"f7",
X"ad",
X"42",
X"02",
X"85",
X"04",
X"ad",
X"43",
X"02",
X"85",
X"05",
X"ad",
X"04",
X"04",
X"85",
X"0c",
X"ad",
X"05",
X"04",
X"85",
X"0d",
X"a0",
X"7f",
X"b9",
X"00",
X"04",
X"91",
X"04",
X"88",
X"10",
X"f8",
X"18",
X"a5",
X"04",
X"69",
X"80",
X"85",
X"04",
X"a5",
X"05",
X"69",
X"00",
X"85",
X"05",
X"ce",
X"41",
X"02",
X"f0",
X"12",
X"ee",
X"0a",
X"03",
X"20",
X"59",
X"c6",
X"10",
X"dc",
X"20",
X"3e",
X"c6",
X"ad",
X"ea",
X"03",
X"d0",
X"ac",
X"f0",
X"f1",
X"ad",
X"ea",
X"03",
X"f0",
X"03",
X"20",
X"59",
X"c6",
X"20",
X"29",
X"c6",
X"b0",
X"9d",
X"20",
X"3b",
X"c6",
X"e6",
X"09",
X"60",
X"18",
X"ad",
X"42",
X"02",
X"69",
X"06",
X"85",
X"04",
X"ad",
X"43",
X"02",
X"69",
X"00",
X"85",
X"05",
X"6c",
X"04",
X"00",
X"6c",
X"0c",
X"00",
X"a2",
X"3d",
X"a0",
X"c4",
X"8a",
X"a2",
X"00",
X"9d",
X"44",
X"03",
X"98",
X"9d",
X"45",
X"03",
X"a9",
X"09",
X"9d",
X"42",
X"03",
X"a9",
X"ff",
X"9d",
X"48",
X"03",
X"4c",
X"56",
X"e4",
X"ad",
X"ea",
X"03",
X"f0",
X"03",
X"4c",
X"7a",
X"e4",
X"a9",
X"52",
X"8d",
X"02",
X"03",
X"a9",
X"01",
X"8d",
X"01",
X"03",
X"4c",
X"53",
X"e4",
X"a5",
X"08",
X"f0",
X"09",
X"a5",
X"09",
X"29",
X"02",
X"f0",
X"27",
X"4c",
X"a0",
X"c6",
X"ad",
X"e9",
X"03",
X"f0",
X"1f",
X"a9",
X"80",
X"85",
X"3e",
X"ee",
X"ea",
X"03",
X"20",
X"7d",
X"e4",
X"20",
X"bb",
X"c5",
X"a9",
X"00",
X"8d",
X"ea",
X"03",
X"8d",
X"e9",
X"03",
X"06",
X"09",
X"a5",
X"0c",
X"85",
X"02",
X"a5",
X"0d",
X"85",
X"03",
X"60",
X"6c",
X"02",
X"00",
X"a9",
X"a0",
X"8d",
X"46",
X"02",
X"a9",
X"80",
X"8d",
X"d5",
X"02",
X"a9",
X"00",
X"8d",
X"d6",
X"02",
X"60",
X"a9",
X"31",
X"8d",
X"00",
X"03",
X"ad",
X"46",
X"02",
X"ae",
X"02",
X"03",
X"e0",
X"21",
X"f0",
X"02",
X"a9",
X"07",
X"8d",
X"06",
X"03",
X"a2",
X"40",
X"ad",
X"02",
X"03",
X"c9",
X"50",
X"f0",
X"04",
X"c9",
X"57",
X"d0",
X"02",
X"a2",
X"80",
X"c9",
X"53",
X"d0",
X"10",
X"a9",
X"ea",
X"8d",
X"04",
X"03",
X"a9",
X"02",
X"8d",
X"05",
X"03",
X"a0",
X"04",
X"a9",
X"00",
X"f0",
X"06",
X"ac",
X"d5",
X"02",
X"ad",
X"d6",
X"02",
X"8e",
X"03",
X"03",
X"8c",
X"08",
X"03",
X"8d",
X"09",
X"03",
X"20",
X"59",
X"e4",
X"10",
X"01",
X"60",
X"ad",
X"02",
X"03",
X"c9",
X"53",
X"d0",
X"0a",
X"20",
X"3a",
X"c7",
X"a0",
X"02",
X"b1",
X"15",
X"8d",
X"46",
X"02",
X"ad",
X"02",
X"03",
X"c9",
X"21",
X"d0",
X"1f",
X"20",
X"3a",
X"c7",
X"a0",
X"fe",
X"c8",
X"c8",
X"b1",
X"15",
X"c9",
X"ff",
X"d0",
X"f8",
X"c8",
X"b1",
X"15",
X"c8",
X"c9",
X"ff",
X"d0",
X"f2",
X"88",
X"88",
X"8c",
X"08",
X"03",
X"a9",
X"00",
X"8d",
X"09",
X"03",
X"ac",
X"03",
X"03",
X"60",
X"ad",
X"04",
X"03",
X"85",
X"15",
X"ad",
X"05",
X"03",
X"85",
X"16",
X"60",
X"a2",
X"05",
X"a9",
X"00",
X"9d",
X"c9",
X"02",
X"ca",
X"10",
X"f8",
X"a9",
X"00",
X"8d",
X"33",
X"02",
X"20",
X"cf",
X"c7",
X"a0",
X"9c",
X"b0",
X"39",
X"8d",
X"88",
X"02",
X"20",
X"cf",
X"c7",
X"a0",
X"9c",
X"b0",
X"2f",
X"8d",
X"45",
X"02",
X"ad",
X"88",
X"02",
X"c9",
X"0b",
X"f0",
X"26",
X"2a",
X"aa",
X"bd",
X"e4",
X"c8",
X"8d",
X"c9",
X"02",
X"bd",
X"e5",
X"c8",
X"8d",
X"ca",
X"02",
X"ad",
X"45",
X"02",
X"cd",
X"33",
X"02",
X"f0",
X"ca",
X"20",
X"cf",
X"c7",
X"a0",
X"9c",
X"b0",
X"08",
X"20",
X"d2",
X"c7",
X"ee",
X"33",
X"02",
X"d0",
X"e9",
X"60",
X"20",
X"cf",
X"c7",
X"a0",
X"9c",
X"b0",
X"2c",
X"8d",
X"c9",
X"02",
X"20",
X"cf",
X"c7",
X"a0",
X"9c",
X"b0",
X"22",
X"8d",
X"ca",
X"02",
X"ad",
X"45",
X"02",
X"c9",
X"01",
X"f0",
X"16",
X"90",
X"17",
X"18",
X"ad",
X"c9",
X"02",
X"6d",
X"d1",
X"02",
X"a8",
X"ad",
X"ca",
X"02",
X"6d",
X"d2",
X"02",
X"8c",
X"c9",
X"02",
X"8d",
X"ca",
X"02",
X"a0",
X"01",
X"60",
X"a0",
X"00",
X"a9",
X"00",
X"f0",
X"f1",
X"6c",
X"cf",
X"02",
X"6c",
X"c9",
X"02",
X"ac",
X"33",
X"02",
X"c0",
X"01",
X"f0",
X"0a",
X"b0",
X"73",
X"8d",
X"4a",
X"02",
X"8d",
X"8e",
X"02",
X"90",
X"6a",
X"8d",
X"4b",
X"02",
X"8d",
X"8f",
X"02",
X"a2",
X"00",
X"ad",
X"88",
X"02",
X"f0",
X"06",
X"c9",
X"0a",
X"f0",
X"15",
X"a2",
X"02",
X"18",
X"ad",
X"4a",
X"02",
X"7d",
X"d1",
X"02",
X"8d",
X"8e",
X"02",
X"ad",
X"4b",
X"02",
X"7d",
X"d2",
X"02",
X"8d",
X"8f",
X"02",
X"18",
X"ad",
X"8e",
X"02",
X"6d",
X"45",
X"02",
X"48",
X"a9",
X"00",
X"6d",
X"8f",
X"02",
X"a8",
X"68",
X"38",
X"e9",
X"02",
X"b0",
X"01",
X"88",
X"48",
X"98",
X"dd",
X"cc",
X"02",
X"68",
X"90",
X"10",
X"d0",
X"05",
X"dd",
X"cb",
X"02",
X"90",
X"09",
X"9d",
X"cb",
X"02",
X"48",
X"98",
X"9d",
X"cc",
X"02",
X"68",
X"ae",
X"88",
X"02",
X"e0",
X"01",
X"f0",
X"10",
X"cc",
X"e6",
X"02",
X"90",
X"0b",
X"d0",
X"05",
X"cd",
X"e5",
X"02",
X"90",
X"04",
X"68",
X"68",
X"a0",
X"9d",
X"60",
X"38",
X"48",
X"ad",
X"33",
X"02",
X"e9",
X"02",
X"18",
X"6d",
X"8e",
X"02",
X"85",
X"36",
X"a9",
X"00",
X"6d",
X"8f",
X"02",
X"85",
X"37",
X"68",
X"a0",
X"00",
X"91",
X"36",
X"4c",
X"50",
X"c8",
X"18",
X"6d",
X"8e",
X"02",
X"85",
X"36",
X"a9",
X"00",
X"6d",
X"8f",
X"02",
X"85",
X"37",
X"a0",
X"00",
X"b1",
X"36",
X"18",
X"6d",
X"d1",
X"02",
X"91",
X"36",
X"e6",
X"36",
X"d0",
X"02",
X"e6",
X"37",
X"b1",
X"36",
X"6d",
X"d2",
X"02",
X"91",
X"36",
X"60",
X"a2",
X"00",
X"ac",
X"88",
X"02",
X"c0",
X"04",
X"90",
X"02",
X"a2",
X"02",
X"18",
X"6d",
X"8e",
X"02",
X"85",
X"36",
X"a9",
X"00",
X"6d",
X"8f",
X"02",
X"85",
X"37",
X"a0",
X"00",
X"b1",
X"36",
X"18",
X"7d",
X"d1",
X"02",
X"91",
X"36",
X"60",
X"48",
X"ad",
X"33",
X"02",
X"6a",
X"68",
X"b0",
X"15",
X"18",
X"6d",
X"8e",
X"02",
X"85",
X"36",
X"a9",
X"00",
X"6d",
X"8f",
X"02",
X"85",
X"37",
X"a0",
X"00",
X"b1",
X"36",
X"8d",
X"88",
X"02",
X"60",
X"18",
X"6d",
X"d1",
X"02",
X"a9",
X"00",
X"6d",
X"d2",
X"02",
X"6d",
X"88",
X"02",
X"a0",
X"00",
X"91",
X"36",
X"f0",
X"ed",
X"d5",
X"c7",
X"d5",
X"c7",
X"92",
X"c8",
X"92",
X"c8",
X"92",
X"c8",
X"92",
X"c8",
X"6d",
X"c8",
X"6d",
X"c8",
X"b5",
X"c8",
X"b5",
X"c8",
X"d5",
X"c7",
X"95",
X"c7",
X"a9",
X"ff",
X"8d",
X"44",
X"02",
X"ad",
X"01",
X"d3",
X"29",
X"7f",
X"8d",
X"01",
X"d3",
X"4c",
X"83",
X"e4",
X"a9",
X"01",
X"8d",
X"48",
X"02",
X"ad",
X"48",
X"02",
X"8d",
X"ff",
X"d1",
X"ad",
X"03",
X"d8",
X"c9",
X"80",
X"d0",
X"0a",
X"ad",
X"0b",
X"d8",
X"c9",
X"91",
X"d0",
X"03",
X"20",
X"19",
X"d8",
X"0e",
X"48",
X"02",
X"d0",
X"e4",
X"a9",
X"00",
X"8d",
X"ff",
X"d1",
X"60",
X"a9",
X"01",
X"8d",
X"42",
X"00",
X"ad",
X"01",
X"03",
X"48",
X"ad",
X"47",
X"02",
X"f0",
X"1a",
X"a2",
X"08",
X"20",
X"af",
X"c9",
X"f0",
X"13",
X"8a",
X"48",
X"20",
X"05",
X"d8",
X"68",
X"aa",
X"90",
X"f2",
X"a9",
X"00",
X"8d",
X"48",
X"02",
X"8d",
X"ff",
X"d1",
X"f0",
X"03",
X"20",
X"71",
X"e9",
X"68",
X"8d",
X"01",
X"03",
X"a9",
X"00",
X"8d",
X"42",
X"00",
X"8c",
X"03",
X"03",
X"ac",
X"03",
X"03",
X"60",
X"a2",
X"08",
X"6a",
X"b0",
X"03",
X"ca",
X"d0",
X"fa",
X"ad",
X"48",
X"02",
X"48",
X"bd",
X"20",
X"ca",
X"8d",
X"48",
X"02",
X"8d",
X"ff",
X"d1",
X"20",
X"08",
X"d8",
X"68",
X"8d",
X"48",
X"02",
X"8d",
X"ff",
X"d1",
X"68",
X"aa",
X"68",
X"40",
X"a0",
X"01",
X"4c",
X"dc",
X"c9",
X"a0",
X"03",
X"4c",
X"dc",
X"c9",
X"a0",
X"05",
X"4c",
X"dc",
X"c9",
X"a0",
X"07",
X"4c",
X"dc",
X"c9",
X"a0",
X"09",
X"4c",
X"dc",
X"c9",
X"a0",
X"0b",
X"4c",
X"dc",
X"c9",
X"ca",
X"10",
X"09",
X"a9",
X"00",
X"8d",
X"48",
X"02",
X"8d",
X"ff",
X"d1",
X"60",
X"ad",
X"47",
X"02",
X"3d",
X"21",
X"ca",
X"f0",
X"ec",
X"8d",
X"48",
X"02",
X"8d",
X"ff",
X"d1",
X"60",
X"b9",
X"0d",
X"d8",
X"48",
X"88",
X"b9",
X"0d",
X"d8",
X"48",
X"ad",
X"4c",
X"02",
X"ae",
X"4d",
X"02",
X"a0",
X"92",
X"60",
X"8d",
X"4c",
X"02",
X"8e",
X"4d",
X"02",
X"ad",
X"42",
X"00",
X"48",
X"a9",
X"01",
X"8d",
X"42",
X"00",
X"a2",
X"08",
X"20",
X"af",
X"c9",
X"f0",
X"11",
X"8a",
X"48",
X"98",
X"48",
X"20",
X"ca",
X"c9",
X"90",
X"20",
X"8d",
X"4c",
X"02",
X"68",
X"68",
X"4c",
X"05",
X"ca",
X"a0",
X"82",
X"a9",
X"00",
X"8d",
X"48",
X"02",
X"8d",
X"ff",
X"d1",
X"68",
X"8d",
X"42",
X"00",
X"ad",
X"4c",
X"02",
X"8c",
X"4d",
X"02",
X"ac",
X"4d",
X"02",
X"60",
X"68",
X"a8",
X"68",
X"aa",
X"90",
X"cc",
X"80",
X"40",
X"20",
X"10",
X"08",
X"04",
X"02",
X"01",
X"ae",
X"2e",
X"00",
X"bd",
X"4d",
X"03",
X"20",
X"de",
X"e7",
X"b0",
X"20",
X"18",
X"20",
X"9e",
X"e8",
X"b0",
X"1a",
X"ae",
X"2e",
X"00",
X"bd",
X"4c",
X"03",
X"20",
X"16",
X"e7",
X"b0",
X"0f",
X"ae",
X"2e",
X"00",
X"9d",
X"40",
X"03",
X"85",
X"20",
X"a9",
X"03",
X"85",
X"17",
X"4c",
X"5c",
X"e5",
X"4c",
X"10",
X"e5",
X"00",
X"13",
X"16",
X"d1",
X"e4",
X"e4",
X"e8",
X"29",
X"eb",
X"ee",
X"00",
X"00",
X"2d",
X"25",
X"2d",
X"2f",
X"32",
X"39",
X"00",
X"34",
X"25",
X"33",
X"34",
X"00",
X"00",
X"00",
X"32",
X"2f",
X"2d",
X"32",
X"21",
X"2d",
X"00",
X"00",
X"2b",
X"25",
X"39",
X"22",
X"2f",
X"21",
X"32",
X"24",
X"00",
X"34",
X"25",
X"33",
X"34",
X"00",
X"00",
X"00",
X"b2",
X"91",
X"00",
X"92",
X"00",
X"93",
X"00",
X"94",
X"00",
X"a8",
X"00",
X"a1",
X"00",
X"a2",
X"00",
X"00",
X"00",
X"5b",
X"00",
X"11",
X"00",
X"12",
X"00",
X"13",
X"00",
X"14",
X"00",
X"15",
X"00",
X"16",
X"00",
X"17",
X"00",
X"18",
X"00",
X"19",
X"00",
X"10",
X"00",
X"1c",
X"00",
X"1e",
X"00",
X"a2",
X"80",
X"b3",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"00",
X"31",
X"00",
X"37",
X"00",
X"25",
X"00",
X"32",
X"00",
X"34",
X"00",
X"39",
X"00",
X"35",
X"00",
X"29",
X"00",
X"2f",
X"00",
X"30",
X"00",
X"0d",
X"00",
X"1d",
X"00",
X"b2",
X"b4",
X"00",
X"00",
X"00",
X"80",
X"dc",
X"80",
X"00",
X"21",
X"00",
X"33",
X"00",
X"24",
X"00",
X"26",
X"00",
X"27",
X"00",
X"28",
X"00",
X"2a",
X"00",
X"2b",
X"00",
X"2c",
X"00",
X"1b",
X"00",
X"0b",
X"00",
X"0a",
X"00",
X"a3",
X"00",
X"00",
X"00",
X"80",
X"b3",
X"a8",
X"80",
X"00",
X"3a",
X"00",
X"38",
X"00",
X"23",
X"00",
X"36",
X"00",
X"22",
X"00",
X"2e",
X"00",
X"2d",
X"00",
X"0c",
X"00",
X"0e",
X"00",
X"0f",
X"00",
X"80",
X"b3",
X"a8",
X"80",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"80",
X"b3",
X"80",
X"b0",
X"80",
X"a1",
X"80",
X"a3",
X"80",
X"a5",
X"80",
X"80",
X"80",
X"a2",
X"80",
X"a1",
X"80",
X"b2",
X"80",
X"00",
X"33",
X"00",
X"30",
X"00",
X"21",
X"00",
X"23",
X"00",
X"25",
X"00",
X"00",
X"00",
X"22",
X"00",
X"21",
X"00",
X"32",
X"00",
X"00",
X"33",
X"28",
X"00",
X"22",
X"00",
X"33",
X"00",
X"5c",
X"00",
X"36",
X"2f",
X"29",
X"23",
X"25",
X"00",
X"03",
X"a0",
X"11",
X"a9",
X"00",
X"18",
X"71",
X"4a",
X"88",
X"10",
X"fb",
X"69",
X"00",
X"49",
X"ff",
X"60",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"18",
X"18",
X"00",
X"18",
X"00",
X"00",
X"66",
X"66",
X"66",
X"00",
X"00",
X"00",
X"00",
X"00",
X"66",
X"ff",
X"66",
X"66",
X"ff",
X"66",
X"00",
X"18",
X"3e",
X"60",
X"3c",
X"06",
X"7c",
X"18",
X"00",
X"00",
X"66",
X"6c",
X"18",
X"30",
X"66",
X"46",
X"00",
X"1c",
X"36",
X"1c",
X"38",
X"6f",
X"66",
X"3b",
X"00",
X"00",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"00",
X"00",
X"0e",
X"1c",
X"18",
X"18",
X"1c",
X"0e",
X"00",
X"00",
X"70",
X"38",
X"18",
X"18",
X"38",
X"70",
X"00",
X"00",
X"66",
X"3c",
X"ff",
X"3c",
X"66",
X"00",
X"00",
X"00",
X"18",
X"18",
X"7e",
X"18",
X"18",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"30",
X"00",
X"00",
X"00",
X"7e",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"00",
X"00",
X"06",
X"0c",
X"18",
X"30",
X"60",
X"40",
X"00",
X"00",
X"3c",
X"66",
X"6e",
X"76",
X"66",
X"3c",
X"00",
X"00",
X"18",
X"38",
X"18",
X"18",
X"18",
X"7e",
X"00",
X"00",
X"3c",
X"66",
X"0c",
X"18",
X"30",
X"7e",
X"00",
X"00",
X"7e",
X"0c",
X"18",
X"0c",
X"66",
X"3c",
X"00",
X"00",
X"0c",
X"1c",
X"3c",
X"6c",
X"7e",
X"0c",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"06",
X"66",
X"3c",
X"00",
X"00",
X"3c",
X"60",
X"7c",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"7e",
X"06",
X"0c",
X"18",
X"30",
X"30",
X"00",
X"00",
X"3c",
X"66",
X"3c",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"3c",
X"66",
X"3e",
X"06",
X"0c",
X"38",
X"00",
X"00",
X"00",
X"18",
X"18",
X"00",
X"18",
X"18",
X"00",
X"00",
X"00",
X"18",
X"18",
X"00",
X"18",
X"18",
X"30",
X"06",
X"0c",
X"18",
X"30",
X"18",
X"0c",
X"06",
X"00",
X"00",
X"00",
X"7e",
X"00",
X"00",
X"7e",
X"00",
X"00",
X"60",
X"30",
X"18",
X"0c",
X"18",
X"30",
X"60",
X"00",
X"00",
X"3c",
X"66",
X"0c",
X"18",
X"00",
X"18",
X"00",
X"00",
X"3c",
X"66",
X"6e",
X"6e",
X"60",
X"3e",
X"00",
X"00",
X"18",
X"3c",
X"66",
X"66",
X"7e",
X"66",
X"00",
X"00",
X"7c",
X"66",
X"7c",
X"66",
X"66",
X"7c",
X"00",
X"00",
X"3c",
X"66",
X"60",
X"60",
X"66",
X"3c",
X"00",
X"00",
X"78",
X"6c",
X"66",
X"66",
X"6c",
X"78",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"60",
X"60",
X"7e",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"60",
X"60",
X"60",
X"00",
X"00",
X"3e",
X"60",
X"60",
X"6e",
X"66",
X"3e",
X"00",
X"00",
X"66",
X"66",
X"7e",
X"66",
X"66",
X"66",
X"00",
X"00",
X"7e",
X"18",
X"18",
X"18",
X"18",
X"7e",
X"00",
X"00",
X"06",
X"06",
X"06",
X"06",
X"66",
X"3c",
X"00",
X"00",
X"66",
X"6c",
X"78",
X"78",
X"6c",
X"66",
X"00",
X"00",
X"60",
X"60",
X"60",
X"60",
X"60",
X"7e",
X"00",
X"00",
X"63",
X"77",
X"7f",
X"6b",
X"63",
X"63",
X"00",
X"00",
X"66",
X"76",
X"7e",
X"7e",
X"6e",
X"66",
X"00",
X"00",
X"3c",
X"66",
X"66",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"7c",
X"60",
X"60",
X"00",
X"00",
X"3c",
X"66",
X"66",
X"66",
X"6c",
X"36",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"7c",
X"6c",
X"66",
X"00",
X"00",
X"3c",
X"60",
X"3c",
X"06",
X"06",
X"3c",
X"00",
X"00",
X"7e",
X"18",
X"18",
X"18",
X"18",
X"18",
X"00",
X"00",
X"66",
X"66",
X"66",
X"66",
X"66",
X"7e",
X"00",
X"00",
X"66",
X"66",
X"66",
X"66",
X"3c",
X"18",
X"00",
X"00",
X"63",
X"63",
X"6b",
X"7f",
X"77",
X"63",
X"00",
X"00",
X"66",
X"66",
X"3c",
X"3c",
X"66",
X"66",
X"00",
X"00",
X"66",
X"66",
X"3c",
X"18",
X"18",
X"18",
X"00",
X"00",
X"7e",
X"0c",
X"18",
X"30",
X"60",
X"7e",
X"00",
X"00",
X"1e",
X"18",
X"18",
X"18",
X"18",
X"1e",
X"00",
X"00",
X"40",
X"60",
X"30",
X"18",
X"0c",
X"06",
X"00",
X"00",
X"78",
X"18",
X"18",
X"18",
X"18",
X"78",
X"00",
X"00",
X"08",
X"1c",
X"36",
X"63",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"00",
X"0c",
X"18",
X"3c",
X"06",
X"3e",
X"66",
X"3e",
X"00",
X"30",
X"18",
X"00",
X"66",
X"66",
X"66",
X"3e",
X"00",
X"36",
X"6c",
X"00",
X"76",
X"76",
X"7e",
X"6e",
X"00",
X"0c",
X"18",
X"7e",
X"60",
X"7c",
X"60",
X"7e",
X"00",
X"00",
X"00",
X"3c",
X"60",
X"60",
X"3c",
X"18",
X"30",
X"3c",
X"66",
X"00",
X"3c",
X"66",
X"66",
X"3c",
X"00",
X"30",
X"18",
X"00",
X"3c",
X"66",
X"66",
X"3c",
X"00",
X"30",
X"18",
X"00",
X"38",
X"18",
X"18",
X"3c",
X"00",
X"1c",
X"30",
X"30",
X"78",
X"30",
X"30",
X"7e",
X"00",
X"00",
X"66",
X"00",
X"38",
X"18",
X"18",
X"3c",
X"00",
X"00",
X"66",
X"00",
X"66",
X"66",
X"66",
X"3e",
X"00",
X"36",
X"00",
X"3c",
X"06",
X"3e",
X"66",
X"3e",
X"00",
X"66",
X"00",
X"3c",
X"66",
X"66",
X"66",
X"3c",
X"00",
X"0c",
X"18",
X"00",
X"66",
X"66",
X"66",
X"3e",
X"00",
X"0c",
X"18",
X"00",
X"3c",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"66",
X"00",
X"3c",
X"66",
X"66",
X"3c",
X"00",
X"66",
X"00",
X"66",
X"66",
X"66",
X"66",
X"7e",
X"00",
X"3c",
X"66",
X"1c",
X"06",
X"3e",
X"66",
X"3e",
X"00",
X"3c",
X"66",
X"00",
X"66",
X"66",
X"66",
X"3e",
X"00",
X"3c",
X"66",
X"00",
X"38",
X"18",
X"18",
X"3c",
X"00",
X"0c",
X"18",
X"3c",
X"66",
X"7e",
X"60",
X"3c",
X"00",
X"30",
X"18",
X"3c",
X"66",
X"7e",
X"60",
X"3c",
X"00",
X"36",
X"6c",
X"00",
X"7c",
X"66",
X"66",
X"66",
X"00",
X"3c",
X"c3",
X"3c",
X"66",
X"7e",
X"60",
X"3c",
X"00",
X"18",
X"00",
X"3c",
X"06",
X"3e",
X"66",
X"3e",
X"00",
X"30",
X"18",
X"3c",
X"06",
X"3e",
X"66",
X"3e",
X"00",
X"18",
X"00",
X"18",
X"3c",
X"66",
X"7e",
X"66",
X"00",
X"78",
X"60",
X"78",
X"60",
X"7e",
X"18",
X"1e",
X"00",
X"00",
X"18",
X"3c",
X"7e",
X"18",
X"18",
X"18",
X"00",
X"00",
X"18",
X"18",
X"18",
X"7e",
X"3c",
X"18",
X"00",
X"00",
X"18",
X"30",
X"7e",
X"30",
X"18",
X"00",
X"00",
X"00",
X"18",
X"0c",
X"7e",
X"0c",
X"18",
X"00",
X"00",
X"18",
X"00",
X"18",
X"18",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"3c",
X"06",
X"3e",
X"66",
X"3e",
X"00",
X"00",
X"60",
X"60",
X"7c",
X"66",
X"66",
X"7c",
X"00",
X"00",
X"00",
X"3c",
X"60",
X"60",
X"60",
X"3c",
X"00",
X"00",
X"06",
X"06",
X"3e",
X"66",
X"66",
X"3e",
X"00",
X"00",
X"00",
X"3c",
X"66",
X"7e",
X"60",
X"3c",
X"00",
X"00",
X"0e",
X"18",
X"3e",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"3e",
X"66",
X"66",
X"3e",
X"06",
X"7c",
X"00",
X"60",
X"60",
X"7c",
X"66",
X"66",
X"66",
X"00",
X"00",
X"18",
X"00",
X"38",
X"18",
X"18",
X"3c",
X"00",
X"00",
X"06",
X"00",
X"06",
X"06",
X"06",
X"06",
X"3c",
X"00",
X"60",
X"60",
X"6c",
X"78",
X"6c",
X"66",
X"00",
X"00",
X"38",
X"18",
X"18",
X"18",
X"18",
X"3c",
X"00",
X"00",
X"00",
X"66",
X"7f",
X"7f",
X"6b",
X"63",
X"00",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"66",
X"66",
X"00",
X"00",
X"00",
X"3c",
X"66",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"7c",
X"60",
X"60",
X"00",
X"00",
X"3e",
X"66",
X"66",
X"3e",
X"06",
X"06",
X"00",
X"00",
X"7c",
X"66",
X"60",
X"60",
X"60",
X"00",
X"00",
X"00",
X"3e",
X"60",
X"3c",
X"06",
X"7c",
X"00",
X"00",
X"18",
X"7e",
X"18",
X"18",
X"18",
X"0e",
X"00",
X"00",
X"00",
X"66",
X"66",
X"66",
X"66",
X"3e",
X"00",
X"00",
X"00",
X"66",
X"66",
X"66",
X"3c",
X"18",
X"00",
X"00",
X"00",
X"63",
X"6b",
X"7f",
X"3e",
X"36",
X"00",
X"00",
X"00",
X"66",
X"3c",
X"18",
X"3c",
X"66",
X"00",
X"00",
X"00",
X"66",
X"66",
X"66",
X"3e",
X"0c",
X"78",
X"00",
X"00",
X"7e",
X"0c",
X"18",
X"30",
X"7e",
X"00",
X"66",
X"66",
X"18",
X"3c",
X"66",
X"7e",
X"66",
X"00",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"00",
X"7e",
X"78",
X"7c",
X"6e",
X"66",
X"06",
X"00",
X"08",
X"18",
X"38",
X"78",
X"38",
X"18",
X"08",
X"00",
X"10",
X"18",
X"1c",
X"1e",
X"1c",
X"18",
X"10",
X"00",
X"4c",
X"09",
X"50",
X"20",
X"86",
X"50",
X"4c",
X"91",
X"52",
X"20",
X"86",
X"50",
X"a9",
X"00",
X"85",
X"80",
X"85",
X"81",
X"85",
X"82",
X"8d",
X"08",
X"d2",
X"a9",
X"03",
X"8d",
X"0f",
X"d2",
X"20",
X"10",
X"55",
X"a9",
X"40",
X"8d",
X"0e",
X"d4",
X"a2",
X"00",
X"20",
X"73",
X"57",
X"a2",
X"3a",
X"a0",
X"51",
X"20",
X"9e",
X"50",
X"a9",
X"d0",
X"8d",
X"00",
X"02",
X"a9",
X"50",
X"8d",
X"01",
X"02",
X"a2",
X"0c",
X"a9",
X"aa",
X"20",
X"2a",
X"57",
X"a2",
X"00",
X"8e",
X"0a",
X"d4",
X"e8",
X"d0",
X"fa",
X"ad",
X"0b",
X"d4",
X"c9",
X"18",
X"b0",
X"f9",
X"a9",
X"10",
X"85",
X"87",
X"a9",
X"c0",
X"8d",
X"0e",
X"d4",
X"ad",
X"1f",
X"d0",
X"29",
X"01",
X"d0",
X"f9",
X"a9",
X"ff",
X"8d",
X"fc",
X"02",
X"a5",
X"86",
X"29",
X"0f",
X"c9",
X"01",
X"f0",
X"10",
X"c9",
X"02",
X"f0",
X"0f",
X"c9",
X"04",
X"f0",
X"0e",
X"a9",
X"88",
X"85",
X"86",
X"a9",
X"ff",
X"85",
X"82",
X"4c",
X"91",
X"52",
X"4c",
X"57",
X"55",
X"4c",
X"50",
X"54",
X"a9",
X"11",
X"85",
X"86",
X"a9",
X"21",
X"8d",
X"2f",
X"02",
X"a9",
X"c0",
X"8d",
X"0e",
X"d4",
X"a9",
X"41",
X"85",
X"83",
X"a9",
X"ff",
X"8d",
X"fc",
X"02",
X"60",
X"85",
X"8a",
X"98",
X"48",
X"8a",
X"48",
X"a9",
X"00",
X"8d",
X"2f",
X"02",
X"8d",
X"dc",
X"02",
X"a9",
X"da",
X"8d",
X"00",
X"02",
X"a9",
X"53",
X"8d",
X"01",
X"02",
X"a2",
X"00",
X"8a",
X"20",
X"2a",
X"57",
X"68",
X"aa",
X"68",
X"a8",
X"8e",
X"30",
X"02",
X"86",
X"84",
X"8c",
X"31",
X"02",
X"84",
X"85",
X"a9",
X"21",
X"8d",
X"2f",
X"02",
X"60",
X"48",
X"8a",
X"48",
X"a2",
X"7a",
X"a5",
X"87",
X"c9",
X"01",
X"f0",
X"1f",
X"29",
X"01",
X"f0",
X"0a",
X"e6",
X"a2",
X"a5",
X"a2",
X"29",
X"20",
X"f0",
X"02",
X"a2",
X"2c",
X"8e",
X"0a",
X"d4",
X"8e",
X"16",
X"d0",
X"18",
X"66",
X"87",
X"a9",
X"00",
X"85",
X"4d",
X"68",
X"aa",
X"68",
X"40",
X"a5",
X"88",
X"d0",
X"16",
X"ad",
X"1f",
X"d0",
X"29",
X"02",
X"d0",
X"1a",
X"a5",
X"86",
X"2a",
X"26",
X"86",
X"a9",
X"20",
X"85",
X"a2",
X"a9",
X"ff",
X"85",
X"88",
X"d0",
X"0b",
X"ad",
X"1f",
X"d0",
X"29",
X"02",
X"f0",
X"04",
X"a9",
X"00",
X"85",
X"88",
X"a5",
X"86",
X"29",
X"0f",
X"09",
X"10",
X"85",
X"87",
X"e6",
X"80",
X"d0",
X"02",
X"e6",
X"81",
X"a5",
X"81",
X"c9",
X"fa",
X"d0",
X"04",
X"58",
X"4c",
X"75",
X"50",
X"4c",
X"d3",
X"50",
X"70",
X"70",
X"70",
X"70",
X"70",
X"47",
X"61",
X"51",
X"70",
X"70",
X"70",
X"4e",
X"00",
X"30",
X"70",
X"f0",
X"c6",
X"71",
X"51",
X"70",
X"86",
X"70",
X"86",
X"70",
X"06",
X"70",
X"70",
X"4e",
X"00",
X"30",
X"70",
X"70",
X"70",
X"42",
X"b1",
X"51",
X"41",
X"3a",
X"51",
X"00",
X"00",
X"00",
X"00",
X"33",
X"25",
X"2c",
X"26",
X"00",
X"34",
X"25",
X"33",
X"34",
X"00",
X"00",
X"00",
X"00",
X"00",
X"2d",
X"25",
X"2d",
X"2f",
X"32",
X"39",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"21",
X"35",
X"24",
X"29",
X"2f",
X"0d",
X"36",
X"29",
X"33",
X"35",
X"21",
X"2c",
X"00",
X"00",
X"00",
X"00",
X"2b",
X"25",
X"39",
X"22",
X"2f",
X"21",
X"32",
X"24",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"21",
X"2c",
X"2c",
X"00",
X"34",
X"25",
X"33",
X"34",
X"33",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"42",
X"b3",
X"a5",
X"ac",
X"a5",
X"a3",
X"b4",
X"56",
X"0c",
X"42",
X"b3",
X"b4",
X"a1",
X"b2",
X"b4",
X"56",
X"2f",
X"32",
X"42",
X"b2",
X"a5",
X"b3",
X"a5",
X"b4",
X"56",
X"00",
X"00",
X"00",
X"70",
X"70",
X"70",
X"46",
X"00",
X"30",
X"70",
X"70",
X"06",
X"70",
X"08",
X"70",
X"70",
X"06",
X"70",
X"08",
X"70",
X"08",
X"70",
X"08",
X"70",
X"08",
X"70",
X"70",
X"70",
X"01",
X"ed",
X"51",
X"a0",
X"40",
X"42",
X"f5",
X"51",
X"01",
X"83",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"42",
X"b2",
X"a5",
X"b3",
X"a5",
X"b4",
X"56",
X"2f",
X"32",
X"42",
X"a8",
X"a5",
X"ac",
X"b0",
X"56",
X"34",
X"2f",
X"00",
X"25",
X"38",
X"29",
X"34",
X"00",
X"00",
X"00",
X"00",
X"00",
X"70",
X"70",
X"70",
X"70",
X"46",
X"00",
X"30",
X"70",
X"70",
X"70",
X"70",
X"02",
X"70",
X"70",
X"02",
X"70",
X"02",
X"70",
X"02",
X"70",
X"02",
X"70",
X"02",
X"70",
X"70",
X"01",
X"ed",
X"51",
X"70",
X"70",
X"70",
X"70",
X"46",
X"71",
X"52",
X"70",
X"06",
X"70",
X"70",
X"4b",
X"00",
X"31",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"0b",
X"70",
X"46",
X"00",
X"30",
X"70",
X"01",
X"ed",
X"51",
X"00",
X"00",
X"21",
X"35",
X"24",
X"29",
X"2f",
X"0d",
X"36",
X"29",
X"33",
X"35",
X"21",
X"2c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"34",
X"25",
X"33",
X"34",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"a2",
X"d1",
X"a0",
X"51",
X"a9",
X"00",
X"20",
X"9e",
X"50",
X"a2",
X"01",
X"20",
X"73",
X"57",
X"a2",
X"00",
X"20",
X"59",
X"57",
X"a2",
X"01",
X"20",
X"59",
X"57",
X"ad",
X"20",
X"30",
X"c9",
X"aa",
X"f0",
X"17",
X"a9",
X"55",
X"20",
X"8e",
X"53",
X"20",
X"b1",
X"53",
X"20",
X"73",
X"ff",
X"b0",
X"05",
X"a9",
X"ff",
X"4c",
X"c4",
X"52",
X"a9",
X"aa",
X"20",
X"8e",
X"53",
X"ad",
X"24",
X"30",
X"c9",
X"aa",
X"f0",
X"17",
X"a9",
X"55",
X"20",
X"99",
X"53",
X"20",
X"b1",
X"53",
X"20",
X"92",
X"ff",
X"b0",
X"05",
X"a9",
X"ff",
X"4c",
X"e2",
X"52",
X"a9",
X"aa",
X"20",
X"99",
X"53",
X"a9",
X"c0",
X"85",
X"8d",
X"a9",
X"04",
X"85",
X"a4",
X"a9",
X"00",
X"85",
X"8e",
X"85",
X"90",
X"85",
X"91",
X"85",
X"8f",
X"a6",
X"8e",
X"bd",
X"38",
X"30",
X"25",
X"8d",
X"c9",
X"80",
X"f0",
X"5c",
X"c9",
X"08",
X"f0",
X"58",
X"a9",
X"44",
X"20",
X"c3",
X"53",
X"a5",
X"a4",
X"20",
X"a4",
X"53",
X"a5",
X"a4",
X"49",
X"0c",
X"85",
X"a4",
X"a2",
X"07",
X"bd",
X"4a",
X"54",
X"c5",
X"91",
X"f0",
X"37",
X"ca",
X"10",
X"f6",
X"a9",
X"04",
X"85",
X"92",
X"a2",
X"00",
X"a0",
X"00",
X"8a",
X"91",
X"90",
X"e8",
X"c8",
X"d0",
X"f9",
X"86",
X"93",
X"a0",
X"00",
X"b1",
X"90",
X"c5",
X"93",
X"d0",
X"10",
X"e6",
X"93",
X"c8",
X"d0",
X"f5",
X"e8",
X"d0",
X"e5",
X"e6",
X"91",
X"c6",
X"92",
X"d0",
X"dd",
X"f0",
X"0e",
X"20",
X"b1",
X"53",
X"a9",
X"88",
X"20",
X"c3",
X"53",
X"4c",
X"5e",
X"53",
X"20",
X"b5",
X"53",
X"a9",
X"cc",
X"20",
X"c3",
X"53",
X"a5",
X"8d",
X"30",
X"26",
X"a9",
X"c0",
X"85",
X"8d",
X"e6",
X"8e",
X"18",
X"a5",
X"8f",
X"69",
X"04",
X"85",
X"91",
X"85",
X"8f",
X"cd",
X"e4",
X"02",
X"d0",
X"81",
X"a5",
X"82",
X"d0",
X"03",
X"4c",
X"a9",
X"52",
X"a9",
X"0c",
X"20",
X"a4",
X"53",
X"20",
X"b5",
X"53",
X"4c",
X"57",
X"55",
X"a9",
X"0c",
X"85",
X"8d",
X"d0",
X"da",
X"a2",
X"04",
X"20",
X"2a",
X"57",
X"29",
X"fc",
X"8d",
X"23",
X"30",
X"60",
X"a2",
X"08",
X"20",
X"2a",
X"57",
X"29",
X"fc",
X"8d",
X"27",
X"30",
X"60",
X"85",
X"a5",
X"ad",
X"01",
X"d3",
X"29",
X"f3",
X"05",
X"a5",
X"8d",
X"01",
X"d3",
X"60",
X"a2",
X"3c",
X"d0",
X"02",
X"a2",
X"96",
X"a0",
X"ff",
X"8c",
X"0a",
X"d4",
X"88",
X"d0",
X"fa",
X"ca",
X"d0",
X"f5",
X"60",
X"48",
X"a6",
X"8e",
X"a5",
X"8d",
X"49",
X"ff",
X"3d",
X"38",
X"30",
X"9d",
X"38",
X"30",
X"68",
X"25",
X"8d",
X"1d",
X"38",
X"30",
X"9d",
X"38",
X"30",
X"60",
X"48",
X"a9",
X"0c",
X"8d",
X"17",
X"d0",
X"ad",
X"c8",
X"02",
X"8d",
X"18",
X"d0",
X"a9",
X"00",
X"85",
X"4d",
X"ad",
X"dc",
X"02",
X"f0",
X"0e",
X"a9",
X"00",
X"8d",
X"dc",
X"02",
X"a9",
X"0c",
X"20",
X"a4",
X"53",
X"58",
X"4c",
X"0c",
X"50",
X"a5",
X"8a",
X"f0",
X"47",
X"ad",
X"1f",
X"d0",
X"29",
X"01",
X"f0",
X"04",
X"a9",
X"b3",
X"d0",
X"02",
X"a9",
X"33",
X"8d",
X"1c",
X"30",
X"ad",
X"1f",
X"d0",
X"29",
X"02",
X"f0",
X"04",
X"a9",
X"f3",
X"d0",
X"02",
X"a9",
X"73",
X"8d",
X"1e",
X"30",
X"ad",
X"1f",
X"d0",
X"29",
X"04",
X"f0",
X"04",
X"a9",
X"af",
X"d0",
X"02",
X"a9",
X"2f",
X"8d",
X"20",
X"30",
X"ad",
X"1f",
X"d0",
X"29",
X"07",
X"c9",
X"07",
X"f0",
X"09",
X"a9",
X"64",
X"8d",
X"02",
X"d2",
X"a9",
X"a8",
X"d0",
X"02",
X"a9",
X"00",
X"8d",
X"03",
X"d2",
X"68",
X"40",
X"00",
X"50",
X"54",
X"30",
X"30",
X"30",
X"a2",
X"00",
X"86",
X"94",
X"a2",
X"03",
X"20",
X"73",
X"57",
X"a2",
X"15",
X"a0",
X"52",
X"a9",
X"ff",
X"20",
X"9e",
X"50",
X"a2",
X"02",
X"20",
X"59",
X"57",
X"a2",
X"07",
X"20",
X"59",
X"57",
X"a5",
X"82",
X"f0",
X"13",
X"a6",
X"94",
X"bd",
X"45",
X"55",
X"e6",
X"94",
X"a6",
X"94",
X"e0",
X"13",
X"d0",
X"14",
X"20",
X"b5",
X"53",
X"4c",
X"91",
X"52",
X"ad",
X"fc",
X"02",
X"c9",
X"ff",
X"f0",
X"f9",
X"c9",
X"c0",
X"b0",
X"f5",
X"ad",
X"fc",
X"02",
X"a2",
X"ff",
X"8e",
X"fc",
X"02",
X"48",
X"29",
X"80",
X"f0",
X"05",
X"a2",
X"08",
X"20",
X"59",
X"57",
X"68",
X"48",
X"29",
X"40",
X"f0",
X"0a",
X"a2",
X"05",
X"20",
X"59",
X"57",
X"a2",
X"04",
X"20",
X"59",
X"57",
X"68",
X"29",
X"3f",
X"c9",
X"21",
X"f0",
X"68",
X"c9",
X"2c",
X"f0",
X"74",
X"c9",
X"34",
X"f0",
X"68",
X"c9",
X"0c",
X"f0",
X"76",
X"aa",
X"bd",
X"9c",
X"57",
X"48",
X"a9",
X"21",
X"85",
X"95",
X"a9",
X"30",
X"85",
X"96",
X"68",
X"a0",
X"ff",
X"c8",
X"d1",
X"95",
X"d0",
X"fb",
X"b1",
X"95",
X"49",
X"80",
X"91",
X"95",
X"a5",
X"82",
X"f0",
X"13",
X"20",
X"05",
X"55",
X"a2",
X"14",
X"20",
X"b7",
X"53",
X"20",
X"10",
X"55",
X"a2",
X"0a",
X"20",
X"b7",
X"53",
X"4c",
X"62",
X"54",
X"20",
X"05",
X"55",
X"ad",
X"0f",
X"d2",
X"29",
X"04",
X"f0",
X"f9",
X"20",
X"10",
X"55",
X"4c",
X"62",
X"54",
X"a9",
X"64",
X"8d",
X"00",
X"d2",
X"a9",
X"a8",
X"8d",
X"01",
X"d2",
X"60",
X"a9",
X"00",
X"8d",
X"01",
X"d2",
X"8d",
X"03",
X"d2",
X"8d",
X"05",
X"d2",
X"8d",
X"07",
X"d2",
X"60",
X"a2",
X"03",
X"20",
X"59",
X"57",
X"4c",
X"de",
X"54",
X"a2",
X"06",
X"20",
X"59",
X"57",
X"4c",
X"de",
X"54",
X"a9",
X"7f",
X"8d",
X"52",
X"30",
X"8d",
X"53",
X"30",
X"d0",
X"a5",
X"a9",
X"32",
X"8d",
X"6d",
X"30",
X"a9",
X"34",
X"8d",
X"6e",
X"30",
X"d0",
X"99",
X"52",
X"08",
X"0a",
X"2b",
X"28",
X"0d",
X"3d",
X"39",
X"2d",
X"1f",
X"30",
X"35",
X"1a",
X"7f",
X"2d",
X"3f",
X"28",
X"0d",
X"a2",
X"02",
X"20",
X"73",
X"57",
X"a9",
X"00",
X"85",
X"97",
X"a9",
X"00",
X"85",
X"98",
X"a2",
X"31",
X"a0",
X"52",
X"a9",
X"00",
X"20",
X"9e",
X"50",
X"a2",
X"09",
X"20",
X"59",
X"57",
X"a5",
X"97",
X"4a",
X"18",
X"69",
X"11",
X"8d",
X"0b",
X"30",
X"a2",
X"0f",
X"a9",
X"ff",
X"9d",
X"50",
X"31",
X"9d",
X"b0",
X"31",
X"9d",
X"10",
X"32",
X"9d",
X"70",
X"32",
X"9d",
X"d0",
X"32",
X"ca",
X"10",
X"ec",
X"a9",
X"00",
X"85",
X"99",
X"a9",
X"0c",
X"85",
X"9a",
X"a6",
X"99",
X"bd",
X"17",
X"57",
X"a8",
X"bd",
X"16",
X"57",
X"aa",
X"a5",
X"9a",
X"20",
X"85",
X"56",
X"18",
X"a5",
X"9a",
X"69",
X"06",
X"85",
X"9a",
X"e6",
X"99",
X"e6",
X"99",
X"a5",
X"99",
X"c9",
X"14",
X"d0",
X"e0",
X"20",
X"b1",
X"53",
X"a2",
X"54",
X"a0",
X"31",
X"a9",
X"00",
X"20",
X"85",
X"56",
X"a9",
X"51",
X"20",
X"6c",
X"56",
X"a2",
X"86",
X"a0",
X"31",
X"a9",
X"00",
X"20",
X"85",
X"56",
X"a9",
X"5b",
X"20",
X"6c",
X"56",
X"a2",
X"f8",
X"a0",
X"30",
X"a9",
X"48",
X"20",
X"85",
X"56",
X"a2",
X"c7",
X"a0",
X"30",
X"a9",
X"54",
X"20",
X"85",
X"56",
X"a2",
X"48",
X"a0",
X"32",
X"a9",
X"4e",
X"20",
X"85",
X"56",
X"a9",
X"44",
X"20",
X"6c",
X"56",
X"a2",
X"ca",
X"a0",
X"30",
X"a9",
X"48",
X"20",
X"85",
X"56",
X"a2",
X"1a",
X"a0",
X"32",
X"a9",
X"4e",
X"20",
X"85",
X"56",
X"a2",
X"ca",
X"a0",
X"31",
X"a9",
X"06",
X"20",
X"85",
X"56",
X"a9",
X"3c",
X"20",
X"6c",
X"56",
X"a2",
X"3c",
X"a0",
X"30",
X"a9",
X"48",
X"20",
X"85",
X"56",
X"a2",
X"8c",
X"a0",
X"31",
X"a9",
X"4e",
X"20",
X"85",
X"56",
X"a2",
X"3c",
X"a0",
X"31",
X"a9",
X"06",
X"20",
X"85",
X"56",
X"a9",
X"2d",
X"20",
X"6c",
X"56",
X"a2",
X"9e",
X"a0",
X"30",
X"a9",
X"48",
X"20",
X"85",
X"56",
X"a2",
X"ee",
X"a0",
X"31",
X"a9",
X"4e",
X"20",
X"85",
X"56",
X"a9",
X"35",
X"20",
X"6c",
X"56",
X"20",
X"b5",
X"53",
X"e6",
X"97",
X"e6",
X"97",
X"a5",
X"97",
X"c9",
X"08",
X"d0",
X"07",
X"a5",
X"82",
X"d0",
X"06",
X"4c",
X"5c",
X"55",
X"4c",
X"60",
X"55",
X"20",
X"b5",
X"53",
X"4c",
X"50",
X"54",
X"a4",
X"97",
X"99",
X"00",
X"d2",
X"a9",
X"a8",
X"99",
X"01",
X"d2",
X"a6",
X"98",
X"bd",
X"b6",
X"56",
X"aa",
X"20",
X"b7",
X"53",
X"e6",
X"98",
X"20",
X"10",
X"55",
X"60",
X"86",
X"9b",
X"84",
X"9c",
X"aa",
X"a0",
X"00",
X"a9",
X"10",
X"85",
X"9d",
X"a9",
X"06",
X"85",
X"a3",
X"bd",
X"bc",
X"56",
X"11",
X"9b",
X"91",
X"9b",
X"20",
X"aa",
X"56",
X"c6",
X"9d",
X"d0",
X"f2",
X"e6",
X"9d",
X"e8",
X"c6",
X"a3",
X"d0",
X"eb",
X"60",
X"18",
X"a5",
X"9b",
X"69",
X"10",
X"85",
X"9b",
X"90",
X"02",
X"e6",
X"9c",
X"60",
X"20",
X"20",
X"20",
X"10",
X"10",
X"20",
X"01",
X"1f",
X"3f",
X"7f",
X"3e",
X"1c",
X"00",
X"41",
X"42",
X"4c",
X"70",
X"40",
X"00",
X"01",
X"02",
X"04",
X"08",
X"10",
X"00",
X"43",
X"44",
X"48",
X"48",
X"48",
X"00",
X"44",
X"22",
X"10",
X"08",
X"07",
X"00",
X"04",
X"08",
X"05",
X"02",
X"00",
X"00",
X"30",
X"48",
X"88",
X"84",
X"84",
X"00",
X"88",
X"88",
X"90",
X"a0",
X"c0",
X"00",
X"f0",
X"88",
X"84",
X"82",
X"82",
X"00",
X"82",
X"82",
X"84",
X"88",
X"f0",
X"00",
X"00",
X"00",
X"00",
X"00",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"00",
X"1c",
X"3e",
X"7f",
X"7e",
X"7c",
X"40",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"04",
X"04",
X"06",
X"05",
X"06",
X"c1",
X"30",
X"21",
X"31",
X"81",
X"31",
X"f1",
X"31",
X"02",
X"30",
X"62",
X"30",
X"22",
X"31",
X"82",
X"31",
X"c2",
X"30",
X"c2",
X"31",
X"48",
X"bd",
X"dc",
X"57",
X"85",
X"9e",
X"bd",
X"dd",
X"57",
X"85",
X"9f",
X"bd",
X"de",
X"57",
X"85",
X"a0",
X"bd",
X"df",
X"57",
X"85",
X"a1",
X"a0",
X"00",
X"68",
X"91",
X"9e",
X"e6",
X"9e",
X"d0",
X"02",
X"e6",
X"9f",
X"48",
X"a5",
X"9e",
X"c5",
X"a0",
X"d0",
X"f0",
X"a5",
X"9f",
X"c5",
X"a1",
X"d0",
X"ea",
X"68",
X"60",
X"bd",
X"57",
X"ca",
X"a8",
X"bd",
X"ec",
X"57",
X"85",
X"9e",
X"bd",
X"f6",
X"57",
X"aa",
X"b9",
X"61",
X"ca",
X"9d",
X"00",
X"30",
X"c8",
X"e8",
X"c6",
X"9e",
X"d0",
X"f4",
X"60",
X"bd",
X"8c",
X"57",
X"8d",
X"c4",
X"02",
X"bd",
X"90",
X"57",
X"8d",
X"c5",
X"02",
X"bd",
X"94",
X"57",
X"8d",
X"c6",
X"02",
X"bd",
X"98",
X"57",
X"8d",
X"c8",
X"02",
X"60",
X"2c",
X"0c",
X"2a",
X"18",
X"0f",
X"32",
X"0c",
X"0e",
X"d2",
X"d6",
X"00",
X"b4",
X"d2",
X"a0",
X"30",
X"b4",
X"2c",
X"2a",
X"1b",
X"91",
X"92",
X"2b",
X"0b",
X"0a",
X"2f",
X"00",
X"30",
X"35",
X"b2",
X"29",
X"0d",
X"1d",
X"36",
X"a8",
X"23",
X"93",
X"94",
X"22",
X"38",
X"3a",
X"14",
X"00",
X"13",
X"16",
X"5b",
X"15",
X"12",
X"11",
X"0c",
X"00",
X"0e",
X"2e",
X"00",
X"2d",
X"0f",
X"a1",
X"32",
X"00",
X"25",
X"39",
X"ff",
X"34",
X"37",
X"31",
X"19",
X"00",
X"10",
X"17",
X"a2",
X"18",
X"1c",
X"1e",
X"26",
X"28",
X"24",
X"00",
X"a3",
X"27",
X"33",
X"21",
X"00",
X"30",
X"ff",
X"3e",
X"20",
X"30",
X"24",
X"30",
X"24",
X"30",
X"28",
X"30",
X"00",
X"30",
X"20",
X"30",
X"13",
X"03",
X"13",
X"13",
X"04",
X"04",
X"03",
X"a8",
X"03",
X"07",
X"00",
X"28",
X"00",
X"b7",
X"92",
X"ab",
X"4c",
X"22",
X"72",
X"04",
X"20",
X"a1",
X"db",
X"20",
X"bb",
X"db",
X"b0",
X"39",
X"a2",
X"ed",
X"a0",
X"04",
X"20",
X"48",
X"da",
X"a2",
X"ff",
X"86",
X"f1",
X"20",
X"44",
X"da",
X"f0",
X"04",
X"a9",
X"ff",
X"85",
X"f0",
X"20",
X"94",
X"db",
X"b0",
X"21",
X"48",
X"a6",
X"d5",
X"d0",
X"11",
X"20",
X"eb",
X"db",
X"68",
X"05",
X"d9",
X"85",
X"d9",
X"a6",
X"f1",
X"30",
X"e6",
X"e8",
X"86",
X"f1",
X"d0",
X"e1",
X"68",
X"a6",
X"f1",
X"10",
X"02",
X"e6",
X"ed",
X"4c",
X"18",
X"d8",
X"60",
X"c9",
X"2e",
X"f0",
X"14",
X"c9",
X"45",
X"f0",
X"19",
X"a6",
X"f0",
X"d0",
X"68",
X"c9",
X"2b",
X"f0",
X"c6",
X"c9",
X"2d",
X"f0",
X"00",
X"85",
X"ee",
X"f0",
X"be",
X"a6",
X"f1",
X"10",
X"58",
X"e8",
X"86",
X"f1",
X"f0",
X"b5",
X"a5",
X"f2",
X"85",
X"ec",
X"20",
X"94",
X"db",
X"b0",
X"37",
X"aa",
X"a5",
X"ed",
X"48",
X"86",
X"ed",
X"20",
X"94",
X"db",
X"b0",
X"17",
X"48",
X"a5",
X"ed",
X"0a",
X"85",
X"ed",
X"0a",
X"0a",
X"65",
X"ed",
X"85",
X"ed",
X"68",
X"18",
X"65",
X"ed",
X"85",
X"ed",
X"a4",
X"f2",
X"20",
X"9d",
X"db",
X"a5",
X"ef",
X"f0",
X"09",
X"a5",
X"ed",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"85",
X"ed",
X"68",
X"18",
X"65",
X"ed",
X"85",
X"ed",
X"d0",
X"13",
X"c9",
X"2b",
X"f0",
X"06",
X"c9",
X"2d",
X"d0",
X"07",
X"85",
X"ef",
X"20",
X"94",
X"db",
X"90",
X"ba",
X"a5",
X"ec",
X"85",
X"f2",
X"c6",
X"f2",
X"a5",
X"ed",
X"a6",
X"f1",
X"30",
X"05",
X"f0",
X"03",
X"38",
X"e5",
X"f1",
X"48",
X"2a",
X"68",
X"6a",
X"85",
X"ed",
X"90",
X"03",
X"20",
X"eb",
X"db",
X"a5",
X"ed",
X"18",
X"69",
X"44",
X"85",
X"d4",
X"20",
X"00",
X"dc",
X"b0",
X"0b",
X"a6",
X"ee",
X"f0",
X"06",
X"a5",
X"d4",
X"09",
X"80",
X"85",
X"d4",
X"18",
X"60",
X"20",
X"51",
X"da",
X"a9",
X"30",
X"8d",
X"7f",
X"05",
X"a5",
X"d4",
X"f0",
X"28",
X"29",
X"7f",
X"c9",
X"3f",
X"90",
X"28",
X"c9",
X"45",
X"b0",
X"24",
X"38",
X"e9",
X"3f",
X"20",
X"70",
X"dc",
X"20",
X"a4",
X"dc",
X"09",
X"80",
X"9d",
X"80",
X"05",
X"ad",
X"80",
X"05",
X"c9",
X"2e",
X"f0",
X"03",
X"4c",
X"88",
X"d9",
X"20",
X"c1",
X"dc",
X"4c",
X"9c",
X"d9",
X"a9",
X"b0",
X"8d",
X"80",
X"05",
X"60",
X"a9",
X"01",
X"20",
X"70",
X"dc",
X"20",
X"a4",
X"dc",
X"e8",
X"86",
X"f2",
X"a5",
X"d4",
X"0a",
X"38",
X"e9",
X"80",
X"ae",
X"80",
X"05",
X"e0",
X"30",
X"f0",
X"17",
X"ae",
X"81",
X"05",
X"ac",
X"82",
X"05",
X"8e",
X"82",
X"05",
X"8c",
X"81",
X"05",
X"a6",
X"f2",
X"e0",
X"02",
X"d0",
X"02",
X"e6",
X"f2",
X"18",
X"69",
X"01",
X"85",
X"ed",
X"a9",
X"45",
X"a4",
X"f2",
X"20",
X"9f",
X"dc",
X"84",
X"f2",
X"a5",
X"ed",
X"10",
X"0b",
X"a9",
X"00",
X"38",
X"e5",
X"ed",
X"85",
X"ed",
X"a9",
X"2d",
X"d0",
X"02",
X"a9",
X"2b",
X"20",
X"9f",
X"dc",
X"a2",
X"00",
X"a5",
X"ed",
X"38",
X"e9",
X"0a",
X"90",
X"03",
X"e8",
X"d0",
X"f8",
X"18",
X"69",
X"0a",
X"48",
X"8a",
X"20",
X"9d",
X"dc",
X"68",
X"09",
X"80",
X"20",
X"9d",
X"dc",
X"ad",
X"80",
X"05",
X"c9",
X"30",
X"d0",
X"0d",
X"18",
X"a5",
X"f3",
X"69",
X"01",
X"85",
X"f3",
X"a5",
X"f4",
X"69",
X"00",
X"85",
X"f4",
X"a5",
X"d4",
X"10",
X"09",
X"20",
X"c1",
X"dc",
X"a0",
X"00",
X"a9",
X"2d",
X"91",
X"f3",
X"60",
X"a5",
X"d4",
X"85",
X"f8",
X"a5",
X"d5",
X"85",
X"f7",
X"20",
X"44",
X"da",
X"f8",
X"a0",
X"10",
X"06",
X"f8",
X"26",
X"f7",
X"a2",
X"03",
X"b5",
X"d4",
X"75",
X"d4",
X"95",
X"d4",
X"ca",
X"d0",
X"f7",
X"88",
X"d0",
X"ee",
X"d8",
X"a9",
X"42",
X"85",
X"d4",
X"4c",
X"00",
X"dc",
X"a9",
X"00",
X"85",
X"f7",
X"85",
X"f8",
X"a5",
X"d4",
X"30",
X"66",
X"c9",
X"43",
X"b0",
X"62",
X"38",
X"e9",
X"40",
X"90",
X"3f",
X"69",
X"00",
X"0a",
X"85",
X"f5",
X"20",
X"5a",
X"da",
X"b0",
X"53",
X"a5",
X"f7",
X"85",
X"f9",
X"a5",
X"f8",
X"85",
X"fa",
X"20",
X"5a",
X"da",
X"b0",
X"46",
X"20",
X"5a",
X"da",
X"b0",
X"41",
X"18",
X"a5",
X"f8",
X"65",
X"fa",
X"85",
X"f8",
X"a5",
X"f7",
X"65",
X"f9",
X"85",
X"f7",
X"b0",
X"32",
X"20",
X"b9",
X"dc",
X"18",
X"65",
X"f8",
X"85",
X"f8",
X"a5",
X"f7",
X"69",
X"00",
X"b0",
X"24",
X"85",
X"f7",
X"c6",
X"f5",
X"d0",
X"c6",
X"20",
X"b9",
X"dc",
X"c9",
X"05",
X"90",
X"0d",
X"18",
X"a5",
X"f8",
X"69",
X"01",
X"85",
X"f8",
X"a5",
X"f7",
X"69",
X"00",
X"85",
X"f7",
X"a5",
X"f8",
X"85",
X"d4",
X"a5",
X"f7",
X"85",
X"d5",
X"18",
X"60",
X"38",
X"60",
X"a2",
X"d4",
X"a0",
X"06",
X"a9",
X"00",
X"95",
X"00",
X"e8",
X"88",
X"d0",
X"fa",
X"60",
X"a9",
X"05",
X"85",
X"f4",
X"a9",
X"80",
X"85",
X"f3",
X"60",
X"18",
X"26",
X"f8",
X"26",
X"f7",
X"60",
X"a5",
X"e0",
X"49",
X"80",
X"85",
X"e0",
X"a5",
X"e0",
X"29",
X"7f",
X"85",
X"f7",
X"a5",
X"d4",
X"29",
X"7f",
X"38",
X"e5",
X"f7",
X"10",
X"10",
X"a2",
X"05",
X"b5",
X"d4",
X"b4",
X"e0",
X"95",
X"e0",
X"98",
X"95",
X"d4",
X"ca",
X"10",
X"f4",
X"30",
X"e1",
X"f0",
X"07",
X"c9",
X"05",
X"b0",
X"19",
X"20",
X"3e",
X"dc",
X"f8",
X"a5",
X"d4",
X"45",
X"e0",
X"30",
X"1e",
X"a2",
X"04",
X"18",
X"b5",
X"d5",
X"75",
X"e1",
X"95",
X"d5",
X"ca",
X"10",
X"f7",
X"d8",
X"b0",
X"03",
X"4c",
X"00",
X"dc",
X"a9",
X"01",
X"20",
X"3a",
X"dc",
X"a9",
X"01",
X"85",
X"d5",
X"4c",
X"00",
X"dc",
X"a2",
X"04",
X"38",
X"b5",
X"d5",
X"f5",
X"e1",
X"95",
X"d5",
X"ca",
X"10",
X"f7",
X"90",
X"04",
X"d8",
X"4c",
X"00",
X"dc",
X"a5",
X"d4",
X"49",
X"80",
X"85",
X"d4",
X"38",
X"a2",
X"04",
X"a9",
X"00",
X"f5",
X"d5",
X"95",
X"d5",
X"ca",
X"10",
X"f7",
X"d8",
X"4c",
X"00",
X"dc",
X"a5",
X"d4",
X"f0",
X"45",
X"a5",
X"e0",
X"f0",
X"3e",
X"20",
X"cf",
X"dc",
X"38",
X"e9",
X"40",
X"38",
X"65",
X"e0",
X"30",
X"38",
X"20",
X"e0",
X"dc",
X"a5",
X"df",
X"29",
X"0f",
X"85",
X"f6",
X"c6",
X"f6",
X"30",
X"06",
X"20",
X"01",
X"dd",
X"4c",
X"f7",
X"da",
X"a5",
X"df",
X"4a",
X"4a",
X"4a",
X"4a",
X"85",
X"f6",
X"c6",
X"f6",
X"30",
X"06",
X"20",
X"05",
X"dd",
X"4c",
X"09",
X"db",
X"20",
X"62",
X"dc",
X"c6",
X"f5",
X"d0",
X"d7",
X"a5",
X"ed",
X"85",
X"d4",
X"4c",
X"04",
X"dc",
X"20",
X"44",
X"da",
X"18",
X"60",
X"38",
X"60",
X"a5",
X"e0",
X"f0",
X"fa",
X"a5",
X"d4",
X"f0",
X"f4",
X"20",
X"cf",
X"dc",
X"38",
X"e5",
X"e0",
X"18",
X"69",
X"40",
X"30",
X"eb",
X"20",
X"e0",
X"dc",
X"e6",
X"f5",
X"4c",
X"4e",
X"db",
X"a2",
X"00",
X"b5",
X"d5",
X"95",
X"d4",
X"e8",
X"e0",
X"0c",
X"d0",
X"f7",
X"a0",
X"05",
X"38",
X"f8",
X"b9",
X"da",
X"00",
X"f9",
X"e6",
X"00",
X"99",
X"da",
X"00",
X"88",
X"10",
X"f4",
X"d8",
X"90",
X"04",
X"e6",
X"d9",
X"d0",
X"e9",
X"20",
X"0f",
X"dd",
X"06",
X"d9",
X"06",
X"d9",
X"06",
X"d9",
X"06",
X"d9",
X"a0",
X"05",
X"38",
X"f8",
X"b9",
X"da",
X"00",
X"f9",
X"e0",
X"00",
X"99",
X"da",
X"00",
X"88",
X"10",
X"f4",
X"d8",
X"90",
X"04",
X"e6",
X"d9",
X"d0",
X"e9",
X"20",
X"09",
X"dd",
X"c6",
X"f5",
X"d0",
X"b5",
X"20",
X"62",
X"dc",
X"4c",
X"1a",
X"db",
X"20",
X"af",
X"db",
X"a4",
X"f2",
X"90",
X"02",
X"b1",
X"f3",
X"c8",
X"84",
X"f2",
X"60",
X"a4",
X"f2",
X"a9",
X"20",
X"d1",
X"f3",
X"d0",
X"03",
X"c8",
X"d0",
X"f9",
X"84",
X"f2",
X"60",
X"a4",
X"f2",
X"b1",
X"f3",
X"38",
X"e9",
X"30",
X"90",
X"18",
X"c9",
X"0a",
X"60",
X"a5",
X"f2",
X"48",
X"20",
X"94",
X"db",
X"90",
X"1f",
X"c9",
X"2e",
X"f0",
X"14",
X"c9",
X"2b",
X"f0",
X"07",
X"c9",
X"2d",
X"f0",
X"03",
X"68",
X"38",
X"60",
X"20",
X"94",
X"db",
X"90",
X"0b",
X"c9",
X"2e",
X"d0",
X"f4",
X"20",
X"94",
X"db",
X"90",
X"02",
X"b0",
X"ed",
X"68",
X"85",
X"f2",
X"18",
X"60",
X"a2",
X"e7",
X"d0",
X"02",
X"a2",
X"d5",
X"a0",
X"04",
X"18",
X"36",
X"04",
X"36",
X"03",
X"36",
X"02",
X"36",
X"01",
X"36",
X"00",
X"26",
X"ec",
X"88",
X"d0",
X"f0",
X"60",
X"a2",
X"00",
X"86",
X"da",
X"a2",
X"04",
X"a5",
X"d4",
X"f0",
X"2e",
X"a5",
X"d5",
X"d0",
X"1a",
X"a0",
X"00",
X"b9",
X"d6",
X"00",
X"99",
X"d5",
X"00",
X"c8",
X"c0",
X"05",
X"90",
X"f5",
X"c6",
X"d4",
X"ca",
X"d0",
X"ea",
X"a5",
X"d5",
X"d0",
X"04",
X"85",
X"d4",
X"18",
X"60",
X"a5",
X"d4",
X"29",
X"7f",
X"c9",
X"71",
X"90",
X"01",
X"60",
X"c9",
X"0f",
X"b0",
X"03",
X"20",
X"44",
X"da",
X"18",
X"60",
X"a2",
X"d4",
X"d0",
X"02",
X"a2",
X"e0",
X"86",
X"f9",
X"85",
X"f7",
X"85",
X"f8",
X"a0",
X"04",
X"b5",
X"04",
X"95",
X"05",
X"ca",
X"88",
X"d0",
X"f8",
X"a9",
X"00",
X"95",
X"05",
X"a6",
X"f9",
X"c6",
X"f7",
X"d0",
X"ec",
X"b5",
X"00",
X"18",
X"65",
X"f8",
X"95",
X"00",
X"60",
X"a2",
X"0a",
X"b5",
X"d4",
X"95",
X"d5",
X"ca",
X"10",
X"f9",
X"a9",
X"00",
X"85",
X"d4",
X"60",
X"85",
X"f7",
X"a2",
X"00",
X"a0",
X"00",
X"20",
X"93",
X"dc",
X"38",
X"e9",
X"01",
X"85",
X"f7",
X"b5",
X"d5",
X"4a",
X"4a",
X"4a",
X"4a",
X"20",
X"9d",
X"dc",
X"b5",
X"d5",
X"29",
X"0f",
X"20",
X"9d",
X"dc",
X"e8",
X"e0",
X"05",
X"90",
X"e3",
X"a5",
X"f7",
X"d0",
X"05",
X"a9",
X"2e",
X"20",
X"9f",
X"dc",
X"60",
X"09",
X"30",
X"99",
X"80",
X"05",
X"c8",
X"60",
X"a2",
X"0a",
X"bd",
X"80",
X"05",
X"c9",
X"2e",
X"f0",
X"07",
X"c9",
X"30",
X"d0",
X"07",
X"ca",
X"d0",
X"f2",
X"ca",
X"bd",
X"80",
X"05",
X"60",
X"20",
X"eb",
X"db",
X"a5",
X"ec",
X"29",
X"0f",
X"60",
X"38",
X"a5",
X"f3",
X"e9",
X"01",
X"85",
X"f3",
X"a5",
X"f4",
X"e9",
X"00",
X"85",
X"f4",
X"60",
X"a5",
X"d4",
X"45",
X"e0",
X"29",
X"80",
X"85",
X"ee",
X"06",
X"e0",
X"46",
X"e0",
X"a5",
X"d4",
X"29",
X"7f",
X"60",
X"05",
X"ee",
X"85",
X"ed",
X"a9",
X"00",
X"85",
X"d4",
X"85",
X"e0",
X"20",
X"28",
X"dd",
X"20",
X"e7",
X"db",
X"a5",
X"ec",
X"29",
X"0f",
X"85",
X"e6",
X"a9",
X"05",
X"85",
X"f5",
X"20",
X"34",
X"dd",
X"20",
X"44",
X"da",
X"60",
X"a2",
X"d9",
X"d0",
X"06",
X"a2",
X"d9",
X"d0",
X"08",
X"a2",
X"df",
X"a0",
X"e5",
X"d0",
X"04",
X"a2",
X"df",
X"a0",
X"eb",
X"a9",
X"05",
X"85",
X"f7",
X"18",
X"f8",
X"b5",
X"00",
X"79",
X"00",
X"00",
X"95",
X"00",
X"ca",
X"88",
X"c6",
X"f7",
X"10",
X"f3",
X"d8",
X"60",
X"a0",
X"05",
X"b9",
X"e0",
X"00",
X"99",
X"e6",
X"00",
X"88",
X"10",
X"f7",
X"60",
X"a0",
X"05",
X"b9",
X"d4",
X"00",
X"99",
X"da",
X"00",
X"88",
X"10",
X"f7",
X"60",
X"86",
X"fe",
X"84",
X"ff",
X"85",
X"ef",
X"a2",
X"e0",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"20",
X"b6",
X"dd",
X"a6",
X"fe",
X"a4",
X"ff",
X"20",
X"89",
X"dd",
X"c6",
X"ef",
X"f0",
X"2d",
X"20",
X"db",
X"da",
X"b0",
X"28",
X"18",
X"a5",
X"fe",
X"69",
X"06",
X"85",
X"fe",
X"90",
X"06",
X"a5",
X"ff",
X"69",
X"00",
X"85",
X"ff",
X"a6",
X"fe",
X"a4",
X"ff",
X"20",
X"98",
X"dd",
X"20",
X"66",
X"da",
X"b0",
X"0d",
X"c6",
X"ef",
X"f0",
X"09",
X"a2",
X"e0",
X"a0",
X"05",
X"20",
X"98",
X"dd",
X"30",
X"d3",
X"60",
X"86",
X"fc",
X"84",
X"fd",
X"a0",
X"05",
X"b1",
X"fc",
X"99",
X"d4",
X"00",
X"88",
X"10",
X"f8",
X"60",
X"86",
X"fc",
X"84",
X"fd",
X"a0",
X"05",
X"b1",
X"fc",
X"99",
X"e0",
X"00",
X"88",
X"10",
X"f8",
X"60",
X"86",
X"fc",
X"84",
X"fd",
X"a0",
X"05",
X"b9",
X"d4",
X"00",
X"91",
X"fc",
X"88",
X"10",
X"f8",
X"60",
X"a2",
X"05",
X"b5",
X"d4",
X"95",
X"e0",
X"ca",
X"10",
X"f9",
X"60",
X"a2",
X"89",
X"a0",
X"de",
X"20",
X"98",
X"dd",
X"20",
X"db",
X"da",
X"b0",
X"7f",
X"a9",
X"00",
X"85",
X"f1",
X"a5",
X"d4",
X"85",
X"f0",
X"29",
X"7f",
X"85",
X"d4",
X"38",
X"e9",
X"40",
X"30",
X"26",
X"c9",
X"04",
X"10",
X"6a",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"20",
X"d2",
X"d9",
X"a5",
X"d4",
X"85",
X"f1",
X"a5",
X"d5",
X"d0",
X"58",
X"20",
X"aa",
X"d9",
X"20",
X"b6",
X"dd",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"89",
X"dd",
X"20",
X"60",
X"da",
X"a9",
X"0a",
X"a2",
X"4d",
X"a0",
X"de",
X"20",
X"40",
X"dd",
X"20",
X"b6",
X"dd",
X"20",
X"db",
X"da",
X"a5",
X"f1",
X"f0",
X"23",
X"18",
X"6a",
X"85",
X"e0",
X"a9",
X"01",
X"90",
X"02",
X"a9",
X"10",
X"85",
X"e1",
X"a2",
X"04",
X"a9",
X"00",
X"95",
X"e2",
X"ca",
X"10",
X"fb",
X"a5",
X"e0",
X"18",
X"69",
X"40",
X"b0",
X"19",
X"30",
X"17",
X"85",
X"e0",
X"20",
X"db",
X"da",
X"a5",
X"f0",
X"10",
X"0d",
X"20",
X"b6",
X"dd",
X"a2",
X"8f",
X"a0",
X"de",
X"20",
X"89",
X"dd",
X"20",
X"28",
X"db",
X"60",
X"38",
X"60",
X"3d",
X"17",
X"94",
X"19",
X"00",
X"00",
X"3d",
X"57",
X"33",
X"05",
X"00",
X"00",
X"3e",
X"05",
X"54",
X"76",
X"62",
X"00",
X"3e",
X"32",
X"19",
X"62",
X"27",
X"00",
X"3f",
X"01",
X"68",
X"60",
X"30",
X"36",
X"3f",
X"07",
X"32",
X"03",
X"27",
X"41",
X"3f",
X"25",
X"43",
X"34",
X"56",
X"75",
X"3f",
X"66",
X"27",
X"37",
X"30",
X"50",
X"40",
X"01",
X"15",
X"12",
X"92",
X"55",
X"3f",
X"99",
X"99",
X"99",
X"99",
X"99",
X"3f",
X"43",
X"42",
X"94",
X"48",
X"19",
X"40",
X"01",
X"00",
X"00",
X"00",
X"00",
X"86",
X"fe",
X"84",
X"ff",
X"a2",
X"e0",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"a6",
X"fe",
X"a4",
X"ff",
X"20",
X"98",
X"dd",
X"20",
X"66",
X"da",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"a2",
X"e0",
X"a0",
X"05",
X"20",
X"89",
X"dd",
X"a6",
X"fe",
X"a4",
X"ff",
X"20",
X"98",
X"dd",
X"20",
X"60",
X"da",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"98",
X"dd",
X"20",
X"28",
X"db",
X"60",
X"a9",
X"01",
X"d0",
X"02",
X"a9",
X"00",
X"85",
X"f0",
X"a5",
X"d4",
X"f0",
X"05",
X"30",
X"03",
X"4c",
X"f6",
X"df",
X"38",
X"60",
X"e9",
X"40",
X"0a",
X"85",
X"f1",
X"a5",
X"d5",
X"29",
X"f0",
X"d0",
X"04",
X"a9",
X"01",
X"d0",
X"04",
X"e6",
X"f1",
X"a9",
X"10",
X"85",
X"e1",
X"a2",
X"04",
X"a9",
X"00",
X"95",
X"e2",
X"ca",
X"10",
X"fb",
X"20",
X"28",
X"db",
X"a2",
X"66",
X"a0",
X"df",
X"20",
X"95",
X"de",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"20",
X"b6",
X"dd",
X"20",
X"db",
X"da",
X"a9",
X"0a",
X"a2",
X"72",
X"a0",
X"df",
X"20",
X"40",
X"dd",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"98",
X"dd",
X"20",
X"db",
X"da",
X"a2",
X"6c",
X"a0",
X"df",
X"20",
X"98",
X"dd",
X"20",
X"66",
X"da",
X"20",
X"b6",
X"dd",
X"a9",
X"00",
X"85",
X"d5",
X"a5",
X"f1",
X"85",
X"d4",
X"10",
X"07",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"85",
X"d4",
X"20",
X"aa",
X"d9",
X"24",
X"f1",
X"10",
X"06",
X"a9",
X"80",
X"05",
X"d4",
X"85",
X"d4",
X"20",
X"66",
X"da",
X"a5",
X"f0",
X"f0",
X"0a",
X"a2",
X"89",
X"a0",
X"de",
X"20",
X"98",
X"dd",
X"20",
X"28",
X"db",
X"18",
X"60",
X"40",
X"03",
X"16",
X"22",
X"77",
X"66",
X"3f",
X"50",
X"00",
X"00",
X"00",
X"00",
X"3f",
X"49",
X"15",
X"57",
X"11",
X"08",
X"bf",
X"51",
X"70",
X"49",
X"47",
X"08",
X"3f",
X"39",
X"20",
X"57",
X"61",
X"95",
X"bf",
X"04",
X"39",
X"63",
X"03",
X"55",
X"3f",
X"10",
X"09",
X"30",
X"12",
X"64",
X"3f",
X"09",
X"39",
X"08",
X"04",
X"60",
X"3f",
X"12",
X"42",
X"58",
X"47",
X"42",
X"3f",
X"17",
X"37",
X"12",
X"06",
X"08",
X"3f",
X"28",
X"95",
X"29",
X"71",
X"17",
X"3f",
X"86",
X"85",
X"88",
X"96",
X"44",
X"3e",
X"16",
X"05",
X"44",
X"49",
X"00",
X"be",
X"95",
X"68",
X"38",
X"45",
X"00",
X"3f",
X"02",
X"68",
X"79",
X"94",
X"16",
X"bf",
X"04",
X"92",
X"78",
X"90",
X"80",
X"3f",
X"07",
X"03",
X"15",
X"20",
X"00",
X"bf",
X"08",
X"92",
X"29",
X"12",
X"44",
X"3f",
X"11",
X"08",
X"40",
X"09",
X"11",
X"bf",
X"14",
X"28",
X"31",
X"56",
X"04",
X"3f",
X"19",
X"99",
X"98",
X"77",
X"44",
X"bf",
X"33",
X"33",
X"33",
X"31",
X"13",
X"3f",
X"99",
X"99",
X"99",
X"99",
X"99",
X"3f",
X"78",
X"53",
X"98",
X"16",
X"34",
X"a5",
X"d4",
X"85",
X"e0",
X"38",
X"4c",
X"e0",
X"de",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"18",
X"18",
X"00",
X"18",
X"00",
X"00",
X"66",
X"66",
X"66",
X"00",
X"00",
X"00",
X"00",
X"00",
X"66",
X"ff",
X"66",
X"66",
X"ff",
X"66",
X"00",
X"18",
X"3e",
X"60",
X"3c",
X"06",
X"7c",
X"18",
X"00",
X"00",
X"66",
X"6c",
X"18",
X"30",
X"66",
X"46",
X"00",
X"1c",
X"36",
X"1c",
X"38",
X"6f",
X"66",
X"3b",
X"00",
X"00",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"00",
X"00",
X"0e",
X"1c",
X"18",
X"18",
X"1c",
X"0e",
X"00",
X"00",
X"70",
X"38",
X"18",
X"18",
X"38",
X"70",
X"00",
X"00",
X"66",
X"3c",
X"ff",
X"3c",
X"66",
X"00",
X"00",
X"00",
X"18",
X"18",
X"7e",
X"18",
X"18",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"30",
X"00",
X"00",
X"00",
X"7e",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"00",
X"00",
X"06",
X"0c",
X"18",
X"30",
X"60",
X"40",
X"00",
X"00",
X"3c",
X"66",
X"6e",
X"76",
X"66",
X"3c",
X"00",
X"00",
X"18",
X"38",
X"18",
X"18",
X"18",
X"7e",
X"00",
X"00",
X"3c",
X"66",
X"0c",
X"18",
X"30",
X"7e",
X"00",
X"00",
X"7e",
X"0c",
X"18",
X"0c",
X"66",
X"3c",
X"00",
X"00",
X"0c",
X"1c",
X"3c",
X"6c",
X"7e",
X"0c",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"06",
X"66",
X"3c",
X"00",
X"00",
X"3c",
X"60",
X"7c",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"7e",
X"06",
X"0c",
X"18",
X"30",
X"30",
X"00",
X"00",
X"3c",
X"66",
X"3c",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"3c",
X"66",
X"3e",
X"06",
X"0c",
X"38",
X"00",
X"00",
X"00",
X"18",
X"18",
X"00",
X"18",
X"18",
X"00",
X"00",
X"00",
X"18",
X"18",
X"00",
X"18",
X"18",
X"30",
X"06",
X"0c",
X"18",
X"30",
X"18",
X"0c",
X"06",
X"00",
X"00",
X"00",
X"7e",
X"00",
X"00",
X"7e",
X"00",
X"00",
X"60",
X"30",
X"18",
X"0c",
X"18",
X"30",
X"60",
X"00",
X"00",
X"3c",
X"66",
X"0c",
X"18",
X"00",
X"18",
X"00",
X"00",
X"3c",
X"66",
X"6e",
X"6e",
X"60",
X"3e",
X"00",
X"00",
X"18",
X"3c",
X"66",
X"66",
X"7e",
X"66",
X"00",
X"00",
X"7c",
X"66",
X"7c",
X"66",
X"66",
X"7c",
X"00",
X"00",
X"3c",
X"66",
X"60",
X"60",
X"66",
X"3c",
X"00",
X"00",
X"78",
X"6c",
X"66",
X"66",
X"6c",
X"78",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"60",
X"60",
X"7e",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"60",
X"60",
X"60",
X"00",
X"00",
X"3e",
X"60",
X"60",
X"6e",
X"66",
X"3e",
X"00",
X"00",
X"66",
X"66",
X"7e",
X"66",
X"66",
X"66",
X"00",
X"00",
X"7e",
X"18",
X"18",
X"18",
X"18",
X"7e",
X"00",
X"00",
X"06",
X"06",
X"06",
X"06",
X"66",
X"3c",
X"00",
X"00",
X"66",
X"6c",
X"78",
X"78",
X"6c",
X"66",
X"00",
X"00",
X"60",
X"60",
X"60",
X"60",
X"60",
X"7e",
X"00",
X"00",
X"63",
X"77",
X"7f",
X"6b",
X"63",
X"63",
X"00",
X"00",
X"66",
X"76",
X"7e",
X"7e",
X"6e",
X"66",
X"00",
X"00",
X"3c",
X"66",
X"66",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"7c",
X"60",
X"60",
X"00",
X"00",
X"3c",
X"66",
X"66",
X"66",
X"6c",
X"36",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"7c",
X"6c",
X"66",
X"00",
X"00",
X"3c",
X"60",
X"3c",
X"06",
X"06",
X"3c",
X"00",
X"00",
X"7e",
X"18",
X"18",
X"18",
X"18",
X"18",
X"00",
X"00",
X"66",
X"66",
X"66",
X"66",
X"66",
X"7e",
X"00",
X"00",
X"66",
X"66",
X"66",
X"66",
X"3c",
X"18",
X"00",
X"00",
X"63",
X"63",
X"6b",
X"7f",
X"77",
X"63",
X"00",
X"00",
X"66",
X"66",
X"3c",
X"3c",
X"66",
X"66",
X"00",
X"00",
X"66",
X"66",
X"3c",
X"18",
X"18",
X"18",
X"00",
X"00",
X"7e",
X"0c",
X"18",
X"30",
X"60",
X"7e",
X"00",
X"00",
X"1e",
X"18",
X"18",
X"18",
X"18",
X"1e",
X"00",
X"00",
X"40",
X"60",
X"30",
X"18",
X"0c",
X"06",
X"00",
X"00",
X"78",
X"18",
X"18",
X"18",
X"18",
X"78",
X"00",
X"00",
X"08",
X"1c",
X"36",
X"63",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"00",
X"00",
X"36",
X"7f",
X"7f",
X"3e",
X"1c",
X"08",
X"00",
X"18",
X"18",
X"18",
X"1f",
X"1f",
X"18",
X"18",
X"18",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"18",
X"18",
X"18",
X"f8",
X"f8",
X"00",
X"00",
X"00",
X"18",
X"18",
X"18",
X"f8",
X"f8",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"f8",
X"f8",
X"18",
X"18",
X"18",
X"03",
X"07",
X"0e",
X"1c",
X"38",
X"70",
X"e0",
X"c0",
X"c0",
X"e0",
X"70",
X"38",
X"1c",
X"0e",
X"07",
X"03",
X"01",
X"03",
X"07",
X"0f",
X"1f",
X"3f",
X"7f",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"0f",
X"0f",
X"0f",
X"0f",
X"80",
X"c0",
X"e0",
X"f0",
X"f8",
X"fc",
X"fe",
X"ff",
X"0f",
X"0f",
X"0f",
X"0f",
X"00",
X"00",
X"00",
X"00",
X"f0",
X"f0",
X"f0",
X"f0",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"f0",
X"f0",
X"f0",
X"f0",
X"00",
X"1c",
X"1c",
X"77",
X"77",
X"08",
X"1c",
X"00",
X"00",
X"00",
X"00",
X"1f",
X"1f",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"18",
X"18",
X"18",
X"ff",
X"ff",
X"18",
X"18",
X"18",
X"00",
X"00",
X"3c",
X"7e",
X"7e",
X"7e",
X"3c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"c0",
X"c0",
X"c0",
X"c0",
X"c0",
X"c0",
X"c0",
X"c0",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"18",
X"18",
X"18",
X"1f",
X"1f",
X"00",
X"00",
X"00",
X"78",
X"60",
X"78",
X"60",
X"7e",
X"18",
X"1e",
X"00",
X"00",
X"18",
X"3c",
X"7e",
X"18",
X"18",
X"18",
X"00",
X"00",
X"18",
X"18",
X"18",
X"7e",
X"3c",
X"18",
X"00",
X"00",
X"18",
X"30",
X"7e",
X"30",
X"18",
X"00",
X"00",
X"00",
X"18",
X"0c",
X"7e",
X"0c",
X"18",
X"00",
X"00",
X"00",
X"18",
X"3c",
X"7e",
X"7e",
X"3c",
X"18",
X"00",
X"00",
X"00",
X"3c",
X"06",
X"3e",
X"66",
X"3e",
X"00",
X"00",
X"60",
X"60",
X"7c",
X"66",
X"66",
X"7c",
X"00",
X"00",
X"00",
X"3c",
X"60",
X"60",
X"60",
X"3c",
X"00",
X"00",
X"06",
X"06",
X"3e",
X"66",
X"66",
X"3e",
X"00",
X"00",
X"00",
X"3c",
X"66",
X"7e",
X"60",
X"3c",
X"00",
X"00",
X"0e",
X"18",
X"3e",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"3e",
X"66",
X"66",
X"3e",
X"06",
X"7c",
X"00",
X"60",
X"60",
X"7c",
X"66",
X"66",
X"66",
X"00",
X"00",
X"18",
X"00",
X"38",
X"18",
X"18",
X"3c",
X"00",
X"00",
X"06",
X"00",
X"06",
X"06",
X"06",
X"06",
X"3c",
X"00",
X"60",
X"60",
X"6c",
X"78",
X"6c",
X"66",
X"00",
X"00",
X"38",
X"18",
X"18",
X"18",
X"18",
X"3c",
X"00",
X"00",
X"00",
X"66",
X"7f",
X"7f",
X"6b",
X"63",
X"00",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"66",
X"66",
X"00",
X"00",
X"00",
X"3c",
X"66",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"7c",
X"60",
X"60",
X"00",
X"00",
X"3e",
X"66",
X"66",
X"3e",
X"06",
X"06",
X"00",
X"00",
X"7c",
X"66",
X"60",
X"60",
X"60",
X"00",
X"00",
X"00",
X"3e",
X"60",
X"3c",
X"06",
X"7c",
X"00",
X"00",
X"18",
X"7e",
X"18",
X"18",
X"18",
X"0e",
X"00",
X"00",
X"00",
X"66",
X"66",
X"66",
X"66",
X"3e",
X"00",
X"00",
X"00",
X"66",
X"66",
X"66",
X"3c",
X"18",
X"00",
X"00",
X"00",
X"63",
X"6b",
X"7f",
X"3e",
X"36",
X"00",
X"00",
X"00",
X"66",
X"3c",
X"18",
X"3c",
X"66",
X"00",
X"00",
X"00",
X"66",
X"66",
X"66",
X"3e",
X"0c",
X"78",
X"00",
X"00",
X"7e",
X"0c",
X"18",
X"30",
X"7e",
X"00",
X"00",
X"18",
X"3c",
X"7e",
X"7e",
X"18",
X"3c",
X"00",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"00",
X"7e",
X"78",
X"7c",
X"6e",
X"66",
X"06",
X"00",
X"08",
X"18",
X"38",
X"78",
X"38",
X"18",
X"08",
X"00",
X"10",
X"18",
X"1c",
X"1e",
X"1c",
X"18",
X"10",
X"00",
X"93",
X"ef",
X"2d",
X"f2",
X"49",
X"f2",
X"af",
X"f2",
X"1d",
X"f2",
X"2c",
X"f2",
X"4c",
X"6e",
X"ef",
X"00",
X"8d",
X"ef",
X"2d",
X"f2",
X"7f",
X"f1",
X"a3",
X"f1",
X"1d",
X"f2",
X"ae",
X"f9",
X"4c",
X"6e",
X"ef",
X"00",
X"1d",
X"f2",
X"1d",
X"f2",
X"fc",
X"f2",
X"2c",
X"f2",
X"1d",
X"f2",
X"2c",
X"f2",
X"4c",
X"6e",
X"ef",
X"00",
X"c1",
X"fe",
X"06",
X"ff",
X"c0",
X"fe",
X"ca",
X"fe",
X"a2",
X"fe",
X"c0",
X"fe",
X"4c",
X"99",
X"fe",
X"00",
X"e5",
X"fc",
X"ce",
X"fd",
X"79",
X"fd",
X"b3",
X"fd",
X"cb",
X"fd",
X"e4",
X"fc",
X"4c",
X"db",
X"fc",
X"00",
X"4c",
X"a3",
X"c6",
X"4c",
X"b3",
X"c6",
X"4c",
X"df",
X"e4",
X"4c",
X"33",
X"c9",
X"4c",
X"72",
X"c2",
X"4c",
X"e2",
X"c0",
X"4c",
X"8a",
X"c2",
X"4c",
X"5c",
X"e9",
X"4c",
X"17",
X"ec",
X"4c",
X"0c",
X"c0",
X"4c",
X"c1",
X"e4",
X"4c",
X"23",
X"f2",
X"4c",
X"90",
X"c2",
X"4c",
X"c8",
X"c2",
X"4c",
X"8d",
X"fd",
X"4c",
X"f7",
X"fc",
X"4c",
X"23",
X"f2",
X"4c",
X"00",
X"50",
X"4c",
X"bc",
X"ee",
X"4c",
X"15",
X"e9",
X"4c",
X"98",
X"e8",
X"90",
X"c9",
X"95",
X"c9",
X"9a",
X"c9",
X"9f",
X"c9",
X"a4",
X"c9",
X"a9",
X"c9",
X"4c",
X"0c",
X"c9",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"60",
X"a2",
X"00",
X"a9",
X"ff",
X"9d",
X"40",
X"03",
X"a9",
X"db",
X"9d",
X"46",
X"03",
X"a9",
X"e4",
X"9d",
X"47",
X"03",
X"8a",
X"18",
X"69",
X"10",
X"aa",
X"c9",
X"80",
X"90",
X"e8",
X"60",
X"a0",
X"85",
X"60",
X"85",
X"2f",
X"86",
X"2e",
X"8a",
X"29",
X"0f",
X"d0",
X"04",
X"e0",
X"80",
X"90",
X"05",
X"a0",
X"86",
X"4c",
X"70",
X"e6",
X"a0",
X"00",
X"bd",
X"40",
X"03",
X"99",
X"20",
X"00",
X"e8",
X"c8",
X"c0",
X"0c",
X"90",
X"f4",
X"a5",
X"20",
X"c9",
X"7f",
X"d0",
X"15",
X"a5",
X"22",
X"c9",
X"0c",
X"f0",
X"71",
X"ad",
X"e9",
X"02",
X"d0",
X"05",
X"a0",
X"82",
X"4c",
X"70",
X"e6",
X"20",
X"29",
X"ca",
X"30",
X"f8",
X"a0",
X"84",
X"a5",
X"22",
X"c9",
X"03",
X"90",
X"25",
X"a8",
X"c0",
X"0e",
X"90",
X"02",
X"a0",
X"0e",
X"84",
X"17",
X"b9",
X"2a",
X"e7",
X"f0",
X"0f",
X"c9",
X"02",
X"f0",
X"48",
X"c9",
X"08",
X"b0",
X"5f",
X"c9",
X"04",
X"f0",
X"76",
X"4c",
X"1e",
X"e6",
X"a5",
X"20",
X"c9",
X"ff",
X"f0",
X"05",
X"a0",
X"81",
X"4c",
X"70",
X"e6",
X"ad",
X"e9",
X"02",
X"d0",
X"27",
X"20",
X"ff",
X"e6",
X"b0",
X"22",
X"a9",
X"00",
X"8d",
X"ea",
X"02",
X"8d",
X"eb",
X"02",
X"20",
X"95",
X"e6",
X"b0",
X"e6",
X"20",
X"ea",
X"e6",
X"a9",
X"0b",
X"85",
X"17",
X"20",
X"95",
X"e6",
X"a5",
X"2c",
X"85",
X"26",
X"a5",
X"2d",
X"85",
X"27",
X"4c",
X"72",
X"e6",
X"20",
X"f9",
X"ee",
X"4c",
X"70",
X"e6",
X"a0",
X"01",
X"84",
X"23",
X"20",
X"95",
X"e6",
X"b0",
X"03",
X"20",
X"ea",
X"e6",
X"a9",
X"ff",
X"85",
X"20",
X"a9",
X"e4",
X"85",
X"27",
X"a9",
X"db",
X"85",
X"26",
X"4c",
X"72",
X"e6",
X"a5",
X"20",
X"c9",
X"ff",
X"d0",
X"05",
X"20",
X"ff",
X"e6",
X"b0",
X"a5",
X"20",
X"95",
X"e6",
X"20",
X"ea",
X"e6",
X"a6",
X"2e",
X"bd",
X"40",
X"03",
X"85",
X"20",
X"4c",
X"72",
X"e6",
X"a5",
X"22",
X"25",
X"2a",
X"d0",
X"05",
X"a0",
X"83",
X"4c",
X"70",
X"e6",
X"20",
X"95",
X"e6",
X"b0",
X"f8",
X"a5",
X"28",
X"05",
X"29",
X"d0",
X"08",
X"20",
X"ea",
X"e6",
X"85",
X"2f",
X"4c",
X"72",
X"e6",
X"20",
X"ea",
X"e6",
X"85",
X"2f",
X"30",
X"41",
X"a0",
X"00",
X"91",
X"24",
X"20",
X"d1",
X"e6",
X"a5",
X"22",
X"29",
X"02",
X"d0",
X"0c",
X"a5",
X"2f",
X"c9",
X"9b",
X"d0",
X"06",
X"20",
X"bb",
X"e6",
X"4c",
X"18",
X"e6",
X"20",
X"bb",
X"e6",
X"d0",
X"db",
X"a5",
X"22",
X"29",
X"02",
X"d0",
X"1d",
X"20",
X"ea",
X"e6",
X"85",
X"2f",
X"30",
X"0a",
X"a5",
X"2f",
X"c9",
X"9b",
X"d0",
X"f3",
X"a9",
X"89",
X"85",
X"23",
X"20",
X"c8",
X"e6",
X"a0",
X"00",
X"a9",
X"9b",
X"91",
X"24",
X"20",
X"d1",
X"e6",
X"20",
X"d8",
X"e6",
X"4c",
X"72",
X"e6",
X"a5",
X"22",
X"25",
X"2a",
X"d0",
X"05",
X"a0",
X"87",
X"4c",
X"70",
X"e6",
X"20",
X"95",
X"e6",
X"b0",
X"f8",
X"a5",
X"28",
X"05",
X"29",
X"d0",
X"06",
X"a5",
X"2f",
X"e6",
X"28",
X"d0",
X"06",
X"a0",
X"00",
X"b1",
X"24",
X"85",
X"2f",
X"20",
X"ea",
X"e6",
X"08",
X"20",
X"d1",
X"e6",
X"20",
X"bb",
X"e6",
X"28",
X"30",
X"1d",
X"a5",
X"22",
X"29",
X"02",
X"d0",
X"06",
X"a5",
X"2f",
X"c9",
X"9b",
X"f0",
X"11",
X"a5",
X"28",
X"05",
X"29",
X"d0",
X"db",
X"a5",
X"22",
X"29",
X"02",
X"d0",
X"05",
X"a9",
X"9b",
X"20",
X"ea",
X"e6",
X"20",
X"d8",
X"e6",
X"4c",
X"72",
X"e6",
X"84",
X"23",
X"a4",
X"2e",
X"b9",
X"44",
X"03",
X"85",
X"24",
X"b9",
X"45",
X"03",
X"85",
X"25",
X"a2",
X"00",
X"8e",
X"e9",
X"02",
X"b5",
X"20",
X"99",
X"40",
X"03",
X"e8",
X"c8",
X"e0",
X"0c",
X"90",
X"f5",
X"a5",
X"2f",
X"a6",
X"2e",
X"a4",
X"23",
X"60",
X"a4",
X"20",
X"c0",
X"22",
X"90",
X"04",
X"a0",
X"85",
X"b0",
X"1b",
X"b9",
X"1b",
X"03",
X"85",
X"2c",
X"b9",
X"1c",
X"03",
X"85",
X"2d",
X"a4",
X"17",
X"b9",
X"2a",
X"e7",
X"a8",
X"b1",
X"2c",
X"aa",
X"c8",
X"b1",
X"2c",
X"85",
X"2d",
X"86",
X"2c",
X"18",
X"60",
X"a5",
X"28",
X"d0",
X"02",
X"c6",
X"29",
X"c6",
X"28",
X"a5",
X"28",
X"05",
X"29",
X"60",
X"a5",
X"24",
X"d0",
X"02",
X"c6",
X"25",
X"c6",
X"24",
X"60",
X"e6",
X"24",
X"d0",
X"02",
X"e6",
X"25",
X"60",
X"a6",
X"2e",
X"38",
X"bd",
X"48",
X"03",
X"e5",
X"28",
X"85",
X"28",
X"bd",
X"49",
X"03",
X"e5",
X"29",
X"85",
X"29",
X"60",
X"a0",
X"92",
X"20",
X"f4",
X"e6",
X"84",
X"23",
X"c0",
X"00",
X"60",
X"aa",
X"a5",
X"2d",
X"48",
X"a5",
X"2c",
X"48",
X"8a",
X"a6",
X"2e",
X"60",
X"38",
X"a0",
X"01",
X"b1",
X"24",
X"e9",
X"31",
X"30",
X"04",
X"c9",
X"09",
X"90",
X"02",
X"a9",
X"00",
X"85",
X"21",
X"e6",
X"21",
X"a0",
X"00",
X"b1",
X"24",
X"f0",
X"0c",
X"a0",
X"21",
X"d9",
X"1a",
X"03",
X"f0",
X"09",
X"88",
X"88",
X"88",
X"10",
X"f6",
X"a0",
X"82",
X"38",
X"60",
X"98",
X"85",
X"20",
X"18",
X"60",
X"00",
X"04",
X"04",
X"04",
X"04",
X"06",
X"06",
X"06",
X"06",
X"02",
X"08",
X"0a",
X"a5",
X"08",
X"f0",
X"25",
X"a9",
X"e9",
X"85",
X"4a",
X"a9",
X"03",
X"85",
X"4b",
X"a0",
X"12",
X"18",
X"b1",
X"4a",
X"aa",
X"c8",
X"71",
X"4a",
X"f0",
X"26",
X"b1",
X"4a",
X"85",
X"4b",
X"86",
X"4a",
X"20",
X"56",
X"cb",
X"d0",
X"1b",
X"20",
X"94",
X"e8",
X"b0",
X"16",
X"90",
X"e3",
X"a9",
X"00",
X"8d",
X"fb",
X"03",
X"8d",
X"fc",
X"03",
X"a9",
X"4f",
X"d0",
X"2d",
X"a9",
X"00",
X"a8",
X"20",
X"be",
X"e7",
X"10",
X"01",
X"60",
X"18",
X"ad",
X"e7",
X"02",
X"6d",
X"ea",
X"02",
X"8d",
X"12",
X"03",
X"ad",
X"e8",
X"02",
X"6d",
X"eb",
X"02",
X"8d",
X"13",
X"03",
X"38",
X"ad",
X"e5",
X"02",
X"ed",
X"12",
X"03",
X"ad",
X"e6",
X"02",
X"ed",
X"13",
X"03",
X"b0",
X"09",
X"a9",
X"4e",
X"a8",
X"20",
X"be",
X"e7",
X"4c",
X"6e",
X"e7",
X"ad",
X"ec",
X"02",
X"ae",
X"e7",
X"02",
X"8e",
X"ec",
X"02",
X"ae",
X"e8",
X"02",
X"8e",
X"ed",
X"02",
X"20",
X"de",
X"e7",
X"30",
X"e3",
X"38",
X"20",
X"9e",
X"e8",
X"b0",
X"dd",
X"90",
X"b0",
X"48",
X"a2",
X"09",
X"bd",
X"d4",
X"e7",
X"9d",
X"00",
X"03",
X"ca",
X"10",
X"f7",
X"8c",
X"0b",
X"03",
X"68",
X"8d",
X"0a",
X"03",
X"4c",
X"59",
X"e4",
X"4f",
X"01",
X"40",
X"40",
X"ea",
X"02",
X"1e",
X"00",
X"04",
X"00",
X"8d",
X"13",
X"03",
X"a2",
X"00",
X"8e",
X"12",
X"03",
X"ca",
X"8e",
X"15",
X"03",
X"ad",
X"ec",
X"02",
X"6a",
X"90",
X"08",
X"ee",
X"ec",
X"02",
X"d0",
X"03",
X"ee",
X"ed",
X"02",
X"ad",
X"ec",
X"02",
X"8d",
X"d1",
X"02",
X"ad",
X"ed",
X"02",
X"8d",
X"d2",
X"02",
X"a9",
X"16",
X"8d",
X"cf",
X"02",
X"a9",
X"e8",
X"8d",
X"d0",
X"02",
X"a9",
X"80",
X"8d",
X"d3",
X"02",
X"4c",
X"45",
X"c7",
X"ae",
X"15",
X"03",
X"e8",
X"8e",
X"15",
X"03",
X"f0",
X"08",
X"ae",
X"15",
X"03",
X"bd",
X"7d",
X"03",
X"18",
X"60",
X"a9",
X"80",
X"8d",
X"15",
X"03",
X"20",
X"33",
X"e8",
X"10",
X"ee",
X"38",
X"60",
X"a2",
X"0b",
X"bd",
X"51",
X"e8",
X"9d",
X"00",
X"03",
X"ca",
X"10",
X"f7",
X"ae",
X"12",
X"03",
X"8e",
X"0a",
X"03",
X"e8",
X"8e",
X"12",
X"03",
X"ad",
X"13",
X"03",
X"8d",
X"00",
X"03",
X"4c",
X"59",
X"e4",
X"00",
X"01",
X"26",
X"40",
X"fd",
X"03",
X"1e",
X"00",
X"80",
X"00",
X"00",
X"00",
X"8c",
X"12",
X"03",
X"8d",
X"13",
X"03",
X"a9",
X"e9",
X"85",
X"4a",
X"a9",
X"03",
X"85",
X"4b",
X"a0",
X"12",
X"b1",
X"4a",
X"aa",
X"c8",
X"b1",
X"4a",
X"cd",
X"13",
X"03",
X"d0",
X"07",
X"ec",
X"12",
X"03",
X"d0",
X"02",
X"18",
X"60",
X"c9",
X"00",
X"d0",
X"06",
X"e0",
X"00",
X"d0",
X"02",
X"38",
X"60",
X"86",
X"4a",
X"85",
X"4b",
X"20",
X"56",
X"cb",
X"d0",
X"f5",
X"f0",
X"d7",
X"38",
X"08",
X"b0",
X"28",
X"8d",
X"ed",
X"02",
X"8c",
X"ec",
X"02",
X"08",
X"a9",
X"00",
X"a8",
X"20",
X"5d",
X"e8",
X"b0",
X"27",
X"a0",
X"12",
X"ad",
X"ec",
X"02",
X"91",
X"4a",
X"aa",
X"c8",
X"ad",
X"ed",
X"02",
X"91",
X"4a",
X"86",
X"4a",
X"85",
X"4b",
X"a9",
X"00",
X"91",
X"4a",
X"88",
X"91",
X"4a",
X"20",
X"00",
X"e9",
X"90",
X"0c",
X"ad",
X"ed",
X"02",
X"ac",
X"ec",
X"02",
X"20",
X"15",
X"e9",
X"28",
X"38",
X"60",
X"28",
X"b0",
X"09",
X"a9",
X"00",
X"a0",
X"10",
X"91",
X"4a",
X"c8",
X"91",
X"4a",
X"18",
X"a0",
X"10",
X"ad",
X"e7",
X"02",
X"71",
X"4a",
X"8d",
X"e7",
X"02",
X"c8",
X"ad",
X"e8",
X"02",
X"71",
X"4a",
X"8d",
X"e8",
X"02",
X"a0",
X"0f",
X"a9",
X"00",
X"91",
X"4a",
X"20",
X"56",
X"cb",
X"a0",
X"0f",
X"91",
X"4a",
X"18",
X"60",
X"18",
X"a5",
X"4a",
X"69",
X"0c",
X"8d",
X"12",
X"03",
X"a5",
X"4b",
X"69",
X"00",
X"8d",
X"13",
X"03",
X"6c",
X"12",
X"03",
X"4c",
X"72",
X"c2",
X"20",
X"5d",
X"e8",
X"b0",
X"3b",
X"a8",
X"a5",
X"4a",
X"48",
X"a5",
X"4b",
X"48",
X"86",
X"4a",
X"84",
X"4b",
X"ad",
X"44",
X"02",
X"d0",
X"0f",
X"a0",
X"10",
X"18",
X"b1",
X"4a",
X"c8",
X"71",
X"4a",
X"d0",
X"1f",
X"20",
X"56",
X"cb",
X"d0",
X"1a",
X"a0",
X"12",
X"b1",
X"4a",
X"aa",
X"c8",
X"b1",
X"4a",
X"a8",
X"68",
X"85",
X"4b",
X"68",
X"85",
X"4a",
X"98",
X"a0",
X"13",
X"91",
X"4a",
X"88",
X"8a",
X"91",
X"4a",
X"18",
X"60",
X"68",
X"68",
X"38",
X"60",
X"00",
X"00",
X"4c",
X"33",
X"c9",
X"a9",
X"3c",
X"8d",
X"02",
X"d3",
X"a9",
X"3c",
X"8d",
X"03",
X"d3",
X"a9",
X"03",
X"8d",
X"32",
X"02",
X"85",
X"41",
X"8d",
X"0f",
X"d2",
X"60",
X"ba",
X"8e",
X"18",
X"03",
X"a9",
X"01",
X"85",
X"42",
X"ad",
X"00",
X"03",
X"c9",
X"60",
X"d0",
X"03",
X"4c",
X"9d",
X"eb",
X"a9",
X"00",
X"8d",
X"0f",
X"03",
X"a9",
X"01",
X"8d",
X"bd",
X"02",
X"a9",
X"0d",
X"8d",
X"9c",
X"02",
X"a9",
X"28",
X"8d",
X"04",
X"d2",
X"a9",
X"00",
X"8d",
X"06",
X"d2",
X"18",
X"ad",
X"00",
X"03",
X"6d",
X"01",
X"03",
X"69",
X"ff",
X"8d",
X"3a",
X"02",
X"ad",
X"02",
X"03",
X"8d",
X"3b",
X"02",
X"ad",
X"0a",
X"03",
X"8d",
X"3c",
X"02",
X"ad",
X"0b",
X"03",
X"8d",
X"3d",
X"02",
X"18",
X"a9",
X"3a",
X"85",
X"32",
X"69",
X"04",
X"85",
X"34",
X"a9",
X"02",
X"85",
X"33",
X"85",
X"35",
X"a9",
X"34",
X"8d",
X"03",
X"d3",
X"20",
X"af",
X"ec",
X"ad",
X"3f",
X"02",
X"d0",
X"03",
X"98",
X"d0",
X"08",
X"ce",
X"9c",
X"02",
X"10",
X"b4",
X"4c",
X"22",
X"ea",
X"ad",
X"03",
X"03",
X"10",
X"0d",
X"a9",
X"0d",
X"8d",
X"9c",
X"02",
X"20",
X"87",
X"eb",
X"20",
X"af",
X"ec",
X"f0",
X"2f",
X"20",
X"9a",
X"ec",
X"a9",
X"00",
X"8d",
X"3f",
X"02",
X"20",
X"c0",
X"ec",
X"f0",
X"12",
X"2c",
X"03",
X"03",
X"70",
X"07",
X"ad",
X"3f",
X"02",
X"d0",
X"18",
X"f0",
X"1e",
X"20",
X"87",
X"eb",
X"20",
X"fd",
X"ea",
X"ad",
X"3f",
X"02",
X"f0",
X"05",
X"ad",
X"19",
X"03",
X"85",
X"30",
X"a5",
X"30",
X"c9",
X"01",
X"f0",
X"08",
X"ce",
X"bd",
X"02",
X"30",
X"03",
X"4c",
X"8d",
X"e9",
X"20",
X"84",
X"ec",
X"a9",
X"00",
X"85",
X"42",
X"a4",
X"30",
X"8c",
X"03",
X"03",
X"60",
X"a9",
X"00",
X"8d",
X"3f",
X"02",
X"18",
X"a9",
X"3e",
X"85",
X"32",
X"69",
X"01",
X"85",
X"34",
X"a9",
X"02",
X"85",
X"33",
X"85",
X"35",
X"a9",
X"ff",
X"85",
X"3c",
X"20",
X"fd",
X"ea",
X"a0",
X"ff",
X"a5",
X"30",
X"c9",
X"01",
X"d0",
X"19",
X"ad",
X"3e",
X"02",
X"c9",
X"41",
X"f0",
X"21",
X"c9",
X"43",
X"f0",
X"1d",
X"c9",
X"45",
X"d0",
X"06",
X"a9",
X"90",
X"85",
X"30",
X"d0",
X"04",
X"a9",
X"8b",
X"85",
X"30",
X"a5",
X"30",
X"c9",
X"8a",
X"f0",
X"07",
X"a9",
X"ff",
X"8d",
X"3f",
X"02",
X"d0",
X"02",
X"a0",
X"00",
X"a5",
X"30",
X"8d",
X"19",
X"03",
X"60",
X"a9",
X"01",
X"85",
X"30",
X"20",
X"17",
X"ec",
X"a0",
X"00",
X"84",
X"31",
X"84",
X"3b",
X"84",
X"3a",
X"b1",
X"32",
X"8d",
X"0d",
X"d2",
X"85",
X"31",
X"a5",
X"11",
X"d0",
X"03",
X"4c",
X"c7",
X"ed",
X"a5",
X"3a",
X"f0",
X"f5",
X"20",
X"84",
X"ec",
X"60",
X"98",
X"48",
X"e6",
X"32",
X"d0",
X"02",
X"e6",
X"33",
X"a5",
X"32",
X"c5",
X"34",
X"a5",
X"33",
X"e5",
X"35",
X"90",
X"1c",
X"a5",
X"3b",
X"d0",
X"0b",
X"a5",
X"31",
X"8d",
X"0d",
X"d2",
X"a9",
X"ff",
X"85",
X"3b",
X"d0",
X"09",
X"a5",
X"10",
X"09",
X"08",
X"85",
X"10",
X"8d",
X"0e",
X"d2",
X"68",
X"a8",
X"68",
X"40",
X"a0",
X"00",
X"b1",
X"32",
X"8d",
X"0d",
X"d2",
X"18",
X"65",
X"31",
X"69",
X"00",
X"85",
X"31",
X"4c",
X"d7",
X"ea",
X"a5",
X"3b",
X"f0",
X"0b",
X"85",
X"3a",
X"a5",
X"10",
X"29",
X"f7",
X"85",
X"10",
X"8d",
X"0e",
X"d2",
X"68",
X"40",
X"a9",
X"00",
X"ac",
X"0f",
X"03",
X"d0",
X"02",
X"85",
X"31",
X"85",
X"38",
X"85",
X"39",
X"a9",
X"01",
X"85",
X"30",
X"20",
X"40",
X"ec",
X"a9",
X"3c",
X"8d",
X"03",
X"d3",
X"a5",
X"11",
X"d0",
X"03",
X"4c",
X"c7",
X"ed",
X"ad",
X"17",
X"03",
X"f0",
X"05",
X"a5",
X"39",
X"f0",
X"f0",
X"60",
X"a9",
X"8a",
X"85",
X"30",
X"60",
X"98",
X"48",
X"ad",
X"0f",
X"d2",
X"8d",
X"0a",
X"d2",
X"30",
X"04",
X"a0",
X"8c",
X"84",
X"30",
X"29",
X"20",
X"d0",
X"04",
X"a0",
X"8e",
X"84",
X"30",
X"a5",
X"38",
X"f0",
X"13",
X"ad",
X"0d",
X"d2",
X"c5",
X"31",
X"f0",
X"04",
X"a0",
X"8f",
X"84",
X"30",
X"a9",
X"ff",
X"85",
X"39",
X"68",
X"a8",
X"68",
X"40",
X"ad",
X"0d",
X"d2",
X"a0",
X"00",
X"91",
X"32",
X"18",
X"65",
X"31",
X"69",
X"00",
X"85",
X"31",
X"e6",
X"32",
X"d0",
X"02",
X"e6",
X"33",
X"a5",
X"32",
X"c5",
X"34",
X"a5",
X"33",
X"e5",
X"35",
X"90",
X"de",
X"a5",
X"3c",
X"f0",
X"06",
X"a9",
X"00",
X"85",
X"3c",
X"f0",
X"d0",
X"a9",
X"ff",
X"85",
X"38",
X"d0",
X"ce",
X"18",
X"ad",
X"04",
X"03",
X"85",
X"32",
X"6d",
X"08",
X"03",
X"85",
X"34",
X"ad",
X"05",
X"03",
X"85",
X"33",
X"6d",
X"09",
X"03",
X"85",
X"35",
X"60",
X"ad",
X"03",
X"03",
X"10",
X"32",
X"a9",
X"cc",
X"8d",
X"04",
X"d2",
X"a9",
X"05",
X"8d",
X"06",
X"d2",
X"20",
X"17",
X"ec",
X"a6",
X"62",
X"bc",
X"15",
X"ee",
X"ad",
X"0b",
X"03",
X"30",
X"03",
X"bc",
X"11",
X"ee",
X"a2",
X"00",
X"20",
X"e2",
X"ed",
X"a9",
X"34",
X"8d",
X"02",
X"d3",
X"ad",
X"17",
X"03",
X"d0",
X"fb",
X"20",
X"87",
X"eb",
X"20",
X"88",
X"ea",
X"4c",
X"04",
X"ec",
X"a9",
X"ff",
X"8d",
X"0f",
X"03",
X"a6",
X"62",
X"bc",
X"17",
X"ee",
X"ad",
X"0b",
X"03",
X"30",
X"03",
X"bc",
X"13",
X"ee",
X"a2",
X"00",
X"20",
X"e2",
X"ed",
X"a9",
X"34",
X"8d",
X"02",
X"d3",
X"ad",
X"17",
X"03",
X"d0",
X"fb",
X"20",
X"87",
X"eb",
X"20",
X"9a",
X"ec",
X"20",
X"e2",
X"ed",
X"20",
X"3d",
X"ed",
X"20",
X"fd",
X"ea",
X"ad",
X"0b",
X"03",
X"30",
X"05",
X"a9",
X"3c",
X"8d",
X"02",
X"d3",
X"4c",
X"2a",
X"ea",
X"a9",
X"00",
X"8d",
X"17",
X"03",
X"60",
X"a9",
X"07",
X"2d",
X"32",
X"02",
X"09",
X"20",
X"ac",
X"00",
X"03",
X"c0",
X"60",
X"d0",
X"0c",
X"09",
X"08",
X"a0",
X"07",
X"8c",
X"02",
X"d2",
X"a0",
X"05",
X"8c",
X"00",
X"d2",
X"8d",
X"32",
X"02",
X"8d",
X"0f",
X"d2",
X"a9",
X"c7",
X"25",
X"10",
X"09",
X"10",
X"4c",
X"56",
X"ec",
X"a9",
X"07",
X"2d",
X"32",
X"02",
X"09",
X"10",
X"8d",
X"32",
X"02",
X"8d",
X"0f",
X"d2",
X"8d",
X"0a",
X"d2",
X"a9",
X"c7",
X"25",
X"10",
X"09",
X"20",
X"85",
X"10",
X"8d",
X"0e",
X"d2",
X"a9",
X"28",
X"8d",
X"08",
X"d2",
X"a2",
X"06",
X"a9",
X"a8",
X"a4",
X"41",
X"d0",
X"02",
X"a9",
X"a0",
X"9d",
X"01",
X"d2",
X"ca",
X"ca",
X"10",
X"f9",
X"a9",
X"a0",
X"8d",
X"05",
X"d2",
X"ac",
X"00",
X"03",
X"c0",
X"60",
X"f0",
X"06",
X"8d",
X"01",
X"d2",
X"8d",
X"03",
X"d2",
X"60",
X"ea",
X"a9",
X"c7",
X"25",
X"10",
X"85",
X"10",
X"8d",
X"0e",
X"d2",
X"a2",
X"06",
X"a9",
X"00",
X"9d",
X"01",
X"d2",
X"ca",
X"ca",
X"10",
X"f9",
X"60",
X"ad",
X"06",
X"03",
X"6a",
X"6a",
X"a8",
X"29",
X"3f",
X"aa",
X"98",
X"6a",
X"29",
X"c0",
X"a8",
X"60",
X"2c",
X"eb",
X"ad",
X"ea",
X"ec",
X"ea",
X"a2",
X"01",
X"a0",
X"ff",
X"88",
X"d0",
X"fd",
X"ca",
X"d0",
X"f8",
X"20",
X"88",
X"ea",
X"a0",
X"02",
X"a2",
X"00",
X"20",
X"e2",
X"ed",
X"20",
X"37",
X"ea",
X"98",
X"60",
X"8d",
X"10",
X"03",
X"8c",
X"11",
X"03",
X"20",
X"2e",
X"ed",
X"8d",
X"10",
X"03",
X"ad",
X"0c",
X"03",
X"20",
X"2e",
X"ed",
X"8d",
X"0c",
X"03",
X"ad",
X"10",
X"03",
X"38",
X"ed",
X"0c",
X"03",
X"8d",
X"12",
X"03",
X"ad",
X"11",
X"03",
X"38",
X"ed",
X"0d",
X"03",
X"a8",
X"a6",
X"62",
X"a9",
X"00",
X"38",
X"fd",
X"19",
X"ee",
X"18",
X"7d",
X"19",
X"ee",
X"88",
X"10",
X"f9",
X"18",
X"6d",
X"12",
X"03",
X"a8",
X"4a",
X"4a",
X"4a",
X"0a",
X"38",
X"e9",
X"16",
X"aa",
X"98",
X"29",
X"07",
X"a8",
X"a9",
X"f5",
X"18",
X"69",
X"0b",
X"88",
X"10",
X"fa",
X"a0",
X"00",
X"38",
X"e9",
X"07",
X"10",
X"01",
X"88",
X"18",
X"7d",
X"f9",
X"ed",
X"8d",
X"ee",
X"02",
X"98",
X"7d",
X"fa",
X"ed",
X"8d",
X"ef",
X"02",
X"60",
X"c9",
X"7c",
X"30",
X"04",
X"38",
X"e9",
X"7c",
X"60",
X"18",
X"a6",
X"62",
X"7d",
X"1b",
X"ee",
X"60",
X"a5",
X"11",
X"d0",
X"03",
X"4c",
X"c7",
X"ed",
X"78",
X"ad",
X"17",
X"03",
X"d0",
X"02",
X"f0",
X"25",
X"ad",
X"0f",
X"d2",
X"29",
X"10",
X"d0",
X"ea",
X"8d",
X"16",
X"03",
X"ae",
X"0b",
X"d4",
X"a4",
X"14",
X"8e",
X"0c",
X"03",
X"8c",
X"0d",
X"03",
X"a2",
X"01",
X"8e",
X"15",
X"03",
X"a0",
X"0a",
X"a5",
X"11",
X"f0",
X"5b",
X"ad",
X"17",
X"03",
X"d0",
X"04",
X"58",
X"4c",
X"27",
X"eb",
X"ad",
X"0f",
X"d2",
X"29",
X"10",
X"cd",
X"16",
X"03",
X"f0",
X"e9",
X"8d",
X"16",
X"03",
X"88",
X"d0",
X"e3",
X"ce",
X"15",
X"03",
X"30",
X"0c",
X"ad",
X"0b",
X"d4",
X"a4",
X"14",
X"20",
X"c8",
X"ec",
X"a0",
X"09",
X"d0",
X"d2",
X"ad",
X"ee",
X"02",
X"8d",
X"04",
X"d2",
X"ad",
X"ef",
X"02",
X"8d",
X"06",
X"d2",
X"a9",
X"00",
X"8d",
X"0f",
X"d2",
X"ad",
X"32",
X"02",
X"8d",
X"0f",
X"d2",
X"a9",
X"55",
X"91",
X"32",
X"c8",
X"91",
X"32",
X"a9",
X"aa",
X"85",
X"31",
X"18",
X"a5",
X"32",
X"69",
X"02",
X"85",
X"32",
X"a5",
X"33",
X"69",
X"00",
X"85",
X"33",
X"58",
X"60",
X"20",
X"84",
X"ec",
X"a9",
X"3c",
X"8d",
X"02",
X"d3",
X"a9",
X"3c",
X"8d",
X"03",
X"d3",
X"a9",
X"80",
X"85",
X"30",
X"ae",
X"18",
X"03",
X"9a",
X"c6",
X"11",
X"58",
X"4c",
X"2a",
X"ea",
X"a9",
X"11",
X"8d",
X"26",
X"02",
X"a9",
X"ec",
X"8d",
X"27",
X"02",
X"a9",
X"01",
X"78",
X"20",
X"5c",
X"e4",
X"a9",
X"01",
X"8d",
X"17",
X"03",
X"58",
X"60",
X"e8",
X"03",
X"43",
X"04",
X"9e",
X"04",
X"f9",
X"04",
X"54",
X"05",
X"af",
X"05",
X"0a",
X"06",
X"65",
X"06",
X"c0",
X"06",
X"1a",
X"07",
X"75",
X"07",
X"d0",
X"07",
X"b4",
X"96",
X"78",
X"64",
X"0f",
X"0d",
X"0a",
X"08",
X"83",
X"9c",
X"07",
X"20",
X"18",
X"10",
X"0a",
X"0a",
X"10",
X"1c",
X"34",
X"64",
X"c4",
X"c4",
X"c4",
X"c4",
X"1c",
X"10",
X"64",
X"c4",
X"17",
X"17",
X"0b",
X"17",
X"2f",
X"2f",
X"5f",
X"5f",
X"61",
X"61",
X"61",
X"61",
X"17",
X"0b",
X"bf",
X"61",
X"13",
X"13",
X"09",
X"13",
X"27",
X"27",
X"4f",
X"4f",
X"41",
X"41",
X"41",
X"41",
X"13",
X"09",
X"9f",
X"41",
X"02",
X"06",
X"07",
X"08",
X"09",
X"0a",
X"0b",
X"0d",
X"0f",
X"0f",
X"0f",
X"0f",
X"04",
X"05",
X"0c",
X"0e",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"01",
X"01",
X"03",
X"02",
X"02",
X"01",
X"01",
X"02",
X"02",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"03",
X"28",
X"14",
X"14",
X"28",
X"50",
X"50",
X"a0",
X"a0",
X"40",
X"50",
X"50",
X"50",
X"28",
X"28",
X"a0",
X"a0",
X"18",
X"18",
X"0c",
X"18",
X"30",
X"30",
X"60",
X"60",
X"c0",
X"c0",
X"c0",
X"c0",
X"18",
X"0c",
X"c0",
X"c0",
X"00",
X"00",
X"00",
X"02",
X"03",
X"02",
X"03",
X"02",
X"03",
X"01",
X"01",
X"01",
X"00",
X"00",
X"03",
X"02",
X"ff",
X"f0",
X"0f",
X"c0",
X"30",
X"0c",
X"03",
X"80",
X"40",
X"20",
X"10",
X"08",
X"04",
X"02",
X"01",
X"48",
X"98",
X"48",
X"8a",
X"a2",
X"00",
X"dd",
X"1a",
X"03",
X"f0",
X"1e",
X"e8",
X"e8",
X"e8",
X"e0",
X"22",
X"30",
X"f4",
X"a2",
X"00",
X"a8",
X"a9",
X"00",
X"dd",
X"1a",
X"03",
X"f0",
X"13",
X"e8",
X"e8",
X"e8",
X"e0",
X"22",
X"30",
X"f4",
X"68",
X"68",
X"a0",
X"ff",
X"38",
X"60",
X"68",
X"a8",
X"68",
X"e8",
X"38",
X"60",
X"98",
X"9d",
X"1a",
X"03",
X"68",
X"9d",
X"1b",
X"03",
X"68",
X"9d",
X"1c",
X"03",
X"18",
X"60",
X"a0",
X"00",
X"b1",
X"24",
X"a4",
X"21",
X"20",
X"be",
X"e7",
X"10",
X"03",
X"a0",
X"82",
X"60",
X"a9",
X"7f",
X"85",
X"20",
X"a9",
X"25",
X"85",
X"26",
X"a9",
X"ef",
X"85",
X"27",
X"ad",
X"ec",
X"02",
X"ae",
X"2e",
X"00",
X"9d",
X"4d",
X"03",
X"a0",
X"00",
X"b1",
X"24",
X"9d",
X"4c",
X"03",
X"a0",
X"01",
X"60",
X"48",
X"8a",
X"48",
X"29",
X"0f",
X"d0",
X"10",
X"e0",
X"80",
X"10",
X"0c",
X"ad",
X"e9",
X"02",
X"d0",
X"0b",
X"a0",
X"82",
X"68",
X"68",
X"c0",
X"00",
X"60",
X"a0",
X"86",
X"30",
X"f7",
X"8e",
X"2e",
X"00",
X"a0",
X"00",
X"bd",
X"40",
X"03",
X"99",
X"20",
X"00",
X"e8",
X"c8",
X"c0",
X"0c",
X"30",
X"f4",
X"20",
X"29",
X"ca",
X"30",
X"e1",
X"68",
X"aa",
X"68",
X"a8",
X"a5",
X"27",
X"48",
X"a5",
X"26",
X"48",
X"98",
X"a0",
X"92",
X"60",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"4c",
X"05",
X"fd",
X"a9",
X"ff",
X"8d",
X"fc",
X"02",
X"ad",
X"e4",
X"02",
X"85",
X"6a",
X"a9",
X"40",
X"8d",
X"be",
X"02",
X"a9",
X"51",
X"85",
X"79",
X"a9",
X"fb",
X"85",
X"7a",
X"a9",
X"11",
X"85",
X"60",
X"a9",
X"fc",
X"85",
X"61",
X"60",
X"a5",
X"2b",
X"29",
X"0f",
X"d0",
X"08",
X"a5",
X"2a",
X"29",
X"0f",
X"85",
X"2a",
X"a9",
X"00",
X"85",
X"57",
X"c9",
X"10",
X"90",
X"05",
X"a9",
X"91",
X"4c",
X"54",
X"f1",
X"a9",
X"e0",
X"8d",
X"f4",
X"02",
X"a9",
X"cc",
X"8d",
X"6b",
X"02",
X"a9",
X"02",
X"8d",
X"f3",
X"02",
X"8d",
X"2f",
X"02",
X"a9",
X"01",
X"85",
X"4c",
X"a9",
X"c0",
X"05",
X"10",
X"85",
X"10",
X"8d",
X"0e",
X"d2",
X"a9",
X"40",
X"8d",
X"0e",
X"d4",
X"2c",
X"6e",
X"02",
X"10",
X"0c",
X"a9",
X"c4",
X"8d",
X"00",
X"02",
X"a9",
X"fc",
X"8d",
X"01",
X"02",
X"a9",
X"c0",
X"8d",
X"0e",
X"d4",
X"a9",
X"00",
X"8d",
X"93",
X"02",
X"85",
X"64",
X"85",
X"7b",
X"8d",
X"f0",
X"02",
X"a0",
X"0e",
X"a9",
X"01",
X"99",
X"a3",
X"02",
X"88",
X"10",
X"fa",
X"a2",
X"04",
X"bd",
X"08",
X"fb",
X"9d",
X"c4",
X"02",
X"ca",
X"10",
X"f7",
X"a4",
X"6a",
X"88",
X"8c",
X"95",
X"02",
X"a9",
X"60",
X"8d",
X"94",
X"02",
X"a6",
X"57",
X"bd",
X"4d",
X"ee",
X"85",
X"51",
X"a5",
X"6a",
X"85",
X"65",
X"bc",
X"1d",
X"ee",
X"a9",
X"28",
X"20",
X"7a",
X"f5",
X"88",
X"d0",
X"f8",
X"ad",
X"6f",
X"02",
X"29",
X"3f",
X"85",
X"67",
X"a8",
X"e0",
X"08",
X"90",
X"1f",
X"e0",
X"0f",
X"f0",
X"0d",
X"e0",
X"0c",
X"b0",
X"17",
X"8a",
X"6a",
X"6a",
X"6a",
X"29",
X"c0",
X"05",
X"67",
X"a8",
X"a9",
X"10",
X"20",
X"7a",
X"f5",
X"e0",
X"0b",
X"d0",
X"05",
X"a9",
X"06",
X"8d",
X"c8",
X"02",
X"8c",
X"6f",
X"02",
X"a5",
X"64",
X"85",
X"58",
X"a5",
X"65",
X"85",
X"59",
X"ad",
X"0b",
X"d4",
X"c9",
X"7a",
X"d0",
X"f9",
X"20",
X"78",
X"f5",
X"bd",
X"5d",
X"ee",
X"f0",
X"06",
X"a9",
X"ff",
X"85",
X"64",
X"c6",
X"65",
X"20",
X"65",
X"f5",
X"a5",
X"64",
X"85",
X"68",
X"a5",
X"65",
X"85",
X"69",
X"a9",
X"41",
X"20",
X"70",
X"f5",
X"86",
X"66",
X"a9",
X"18",
X"8d",
X"bf",
X"02",
X"a5",
X"57",
X"c9",
X"0c",
X"b0",
X"04",
X"c9",
X"09",
X"b0",
X"39",
X"a5",
X"2a",
X"29",
X"10",
X"f0",
X"33",
X"a9",
X"04",
X"8d",
X"bf",
X"02",
X"a2",
X"02",
X"ad",
X"6e",
X"02",
X"f0",
X"03",
X"20",
X"a0",
X"f5",
X"a9",
X"02",
X"20",
X"69",
X"f5",
X"ca",
X"10",
X"f8",
X"a4",
X"6a",
X"88",
X"98",
X"20",
X"70",
X"f5",
X"a9",
X"60",
X"20",
X"70",
X"f5",
X"a9",
X"42",
X"20",
X"69",
X"f5",
X"18",
X"a9",
X"10",
X"65",
X"66",
X"a8",
X"be",
X"2d",
X"ee",
X"d0",
X"15",
X"a4",
X"66",
X"be",
X"2d",
X"ee",
X"a5",
X"57",
X"d0",
X"0c",
X"ad",
X"6e",
X"02",
X"f0",
X"07",
X"20",
X"a0",
X"f5",
X"a9",
X"22",
X"85",
X"51",
X"a5",
X"51",
X"20",
X"70",
X"f5",
X"ca",
X"d0",
X"f8",
X"a5",
X"57",
X"c9",
X"08",
X"90",
X"26",
X"c9",
X"0f",
X"f0",
X"04",
X"c9",
X"0c",
X"b0",
X"1e",
X"a2",
X"5d",
X"a5",
X"6a",
X"38",
X"e9",
X"10",
X"20",
X"70",
X"f5",
X"a9",
X"00",
X"20",
X"70",
X"f5",
X"a5",
X"51",
X"09",
X"40",
X"20",
X"70",
X"f5",
X"a5",
X"51",
X"20",
X"70",
X"f5",
X"ca",
X"d0",
X"f8",
X"a5",
X"59",
X"20",
X"70",
X"f5",
X"a5",
X"58",
X"20",
X"70",
X"f5",
X"a5",
X"51",
X"09",
X"40",
X"20",
X"70",
X"f5",
X"a9",
X"70",
X"20",
X"70",
X"f5",
X"a9",
X"70",
X"20",
X"70",
X"f5",
X"a5",
X"64",
X"8d",
X"30",
X"02",
X"a5",
X"65",
X"8d",
X"31",
X"02",
X"a9",
X"70",
X"20",
X"70",
X"f5",
X"a5",
X"64",
X"8d",
X"e5",
X"02",
X"a5",
X"65",
X"8d",
X"e6",
X"02",
X"a0",
X"01",
X"ad",
X"30",
X"02",
X"91",
X"68",
X"c8",
X"ad",
X"31",
X"02",
X"91",
X"68",
X"a5",
X"4c",
X"10",
X"10",
X"8d",
X"ec",
X"03",
X"20",
X"94",
X"ef",
X"ad",
X"ec",
X"03",
X"a0",
X"00",
X"8c",
X"ec",
X"03",
X"a8",
X"60",
X"a5",
X"2a",
X"29",
X"20",
X"d0",
X"0b",
X"20",
X"20",
X"f4",
X"8d",
X"90",
X"02",
X"a5",
X"52",
X"8d",
X"91",
X"02",
X"a9",
X"22",
X"0d",
X"2f",
X"02",
X"8d",
X"2f",
X"02",
X"4c",
X"0b",
X"f2",
X"20",
X"ca",
X"f6",
X"20",
X"8f",
X"f1",
X"20",
X"6a",
X"f7",
X"20",
X"0a",
X"f6",
X"4c",
X"1e",
X"f2",
X"20",
X"ac",
X"f5",
X"b1",
X"64",
X"2d",
X"a0",
X"02",
X"46",
X"6f",
X"b0",
X"03",
X"4a",
X"10",
X"f9",
X"8d",
X"fa",
X"02",
X"c9",
X"00",
X"60",
X"8d",
X"fb",
X"02",
X"c9",
X"7d",
X"d0",
X"06",
X"20",
X"20",
X"f4",
X"4c",
X"0b",
X"f2",
X"20",
X"ca",
X"f6",
X"ad",
X"fb",
X"02",
X"c9",
X"9b",
X"d0",
X"06",
X"20",
X"61",
X"f6",
X"4c",
X"0b",
X"f2",
X"20",
X"ca",
X"f1",
X"20",
X"0e",
X"f6",
X"4c",
X"0b",
X"f2",
X"ad",
X"ff",
X"02",
X"d0",
X"fb",
X"a2",
X"02",
X"b5",
X"54",
X"95",
X"5a",
X"ca",
X"10",
X"f9",
X"ad",
X"fb",
X"02",
X"a8",
X"2a",
X"2a",
X"2a",
X"2a",
X"29",
X"03",
X"aa",
X"98",
X"29",
X"9f",
X"1d",
X"49",
X"fb",
X"8d",
X"fa",
X"02",
X"20",
X"ac",
X"f5",
X"ad",
X"fa",
X"02",
X"46",
X"6f",
X"b0",
X"04",
X"0a",
X"4c",
X"f2",
X"f1",
X"2d",
X"a0",
X"02",
X"85",
X"50",
X"ad",
X"a0",
X"02",
X"49",
X"ff",
X"31",
X"64",
X"05",
X"50",
X"91",
X"64",
X"60",
X"20",
X"8f",
X"f1",
X"85",
X"5d",
X"a6",
X"57",
X"d0",
X"0a",
X"ae",
X"f0",
X"02",
X"d0",
X"05",
X"49",
X"80",
X"20",
X"e9",
X"f1",
X"a4",
X"4c",
X"4c",
X"26",
X"f2",
X"4c",
X"fc",
X"c8",
X"a9",
X"01",
X"85",
X"4c",
X"ad",
X"fb",
X"02",
X"60",
X"2c",
X"6e",
X"02",
X"10",
X"eb",
X"a9",
X"40",
X"8d",
X"0e",
X"d4",
X"a9",
X"00",
X"8d",
X"6e",
X"02",
X"a9",
X"ce",
X"8d",
X"00",
X"02",
X"a9",
X"c0",
X"8d",
X"01",
X"02",
X"4c",
X"94",
X"ef",
X"20",
X"62",
X"f9",
X"20",
X"bc",
X"f6",
X"a5",
X"6b",
X"d0",
X"34",
X"a5",
X"54",
X"85",
X"6c",
X"a5",
X"55",
X"85",
X"6d",
X"20",
X"fd",
X"f2",
X"84",
X"4c",
X"ad",
X"fb",
X"02",
X"c9",
X"9b",
X"f0",
X"12",
X"20",
X"be",
X"f2",
X"20",
X"62",
X"f9",
X"a5",
X"63",
X"c9",
X"71",
X"d0",
X"03",
X"20",
X"56",
X"f5",
X"4c",
X"5c",
X"f2",
X"20",
X"18",
X"f7",
X"20",
X"b1",
X"f8",
X"a5",
X"6c",
X"85",
X"54",
X"a5",
X"6d",
X"85",
X"55",
X"a5",
X"6b",
X"f0",
X"11",
X"c6",
X"6b",
X"f0",
X"0d",
X"a5",
X"4c",
X"30",
X"f8",
X"20",
X"80",
X"f1",
X"8d",
X"fb",
X"02",
X"4c",
X"62",
X"f9",
X"20",
X"61",
X"f6",
X"a9",
X"9b",
X"8d",
X"fb",
X"02",
X"20",
X"0b",
X"f2",
X"84",
X"4c",
X"4c",
X"62",
X"f9",
X"6c",
X"64",
X"00",
X"8d",
X"fb",
X"02",
X"20",
X"62",
X"f9",
X"20",
X"bc",
X"f6",
X"a9",
X"00",
X"8d",
X"e8",
X"03",
X"20",
X"18",
X"f7",
X"20",
X"3c",
X"f9",
X"f0",
X"09",
X"0e",
X"a2",
X"02",
X"20",
X"b4",
X"f1",
X"4c",
X"62",
X"f9",
X"ad",
X"fe",
X"02",
X"0d",
X"a2",
X"02",
X"d0",
X"ef",
X"0e",
X"a2",
X"02",
X"e8",
X"ad",
X"e8",
X"03",
X"f0",
X"05",
X"8a",
X"18",
X"69",
X"2d",
X"aa",
X"bd",
X"0d",
X"fb",
X"85",
X"64",
X"bd",
X"0e",
X"fb",
X"85",
X"65",
X"20",
X"ad",
X"f2",
X"20",
X"0b",
X"f2",
X"4c",
X"62",
X"f9",
X"a9",
X"ff",
X"8d",
X"fc",
X"02",
X"a9",
X"00",
X"8d",
X"e8",
X"03",
X"a5",
X"2a",
X"4a",
X"b0",
X"6f",
X"a9",
X"80",
X"a6",
X"11",
X"f0",
X"65",
X"ad",
X"fc",
X"02",
X"c9",
X"ff",
X"f0",
X"e9",
X"85",
X"7c",
X"a2",
X"ff",
X"8e",
X"fc",
X"02",
X"ae",
X"db",
X"02",
X"d0",
X"03",
X"20",
X"83",
X"f9",
X"a8",
X"c0",
X"c0",
X"b0",
X"d0",
X"b1",
X"79",
X"8d",
X"fb",
X"02",
X"aa",
X"30",
X"03",
X"4c",
X"b4",
X"f3",
X"c9",
X"80",
X"f0",
X"c1",
X"c9",
X"81",
X"d0",
X"0a",
X"ad",
X"b6",
X"02",
X"49",
X"80",
X"8d",
X"b6",
X"02",
X"b0",
X"b3",
X"c9",
X"82",
X"d0",
X"0c",
X"ad",
X"be",
X"02",
X"f0",
X"0b",
X"a9",
X"00",
X"8d",
X"be",
X"02",
X"f0",
X"a3",
X"c9",
X"83",
X"d0",
X"07",
X"a9",
X"40",
X"8d",
X"be",
X"02",
X"d0",
X"98",
X"c9",
X"84",
X"d0",
X"08",
X"a9",
X"80",
X"8d",
X"be",
X"02",
X"4c",
X"f8",
X"f2",
X"c9",
X"85",
X"d0",
X"0b",
X"a9",
X"88",
X"85",
X"4c",
X"85",
X"11",
X"a9",
X"9b",
X"4c",
X"da",
X"f3",
X"c9",
X"89",
X"d0",
X"10",
X"ad",
X"db",
X"02",
X"49",
X"ff",
X"8d",
X"db",
X"02",
X"d0",
X"03",
X"20",
X"83",
X"f9",
X"4c",
X"f8",
X"f2",
X"c9",
X"8e",
X"b0",
X"12",
X"c9",
X"8a",
X"90",
X"f5",
X"e9",
X"8a",
X"06",
X"7c",
X"10",
X"02",
X"09",
X"04",
X"a8",
X"b1",
X"60",
X"4c",
X"2a",
X"f3",
X"c9",
X"92",
X"b0",
X"0b",
X"c9",
X"8e",
X"90",
X"df",
X"e9",
X"72",
X"ee",
X"e8",
X"03",
X"d0",
X"26",
X"a5",
X"7c",
X"c9",
X"40",
X"b0",
X"15",
X"ad",
X"fb",
X"02",
X"c9",
X"61",
X"90",
X"0e",
X"c9",
X"7b",
X"b0",
X"0a",
X"ad",
X"be",
X"02",
X"f0",
X"05",
X"05",
X"7c",
X"4c",
X"23",
X"f3",
X"20",
X"3c",
X"f9",
X"f0",
X"09",
X"ad",
X"fb",
X"02",
X"4d",
X"b6",
X"02",
X"8d",
X"fb",
X"02",
X"4c",
X"1e",
X"f2",
X"a9",
X"80",
X"8d",
X"a2",
X"02",
X"60",
X"c6",
X"54",
X"10",
X"06",
X"ae",
X"bf",
X"02",
X"ca",
X"86",
X"54",
X"4c",
X"0c",
X"f9",
X"e6",
X"54",
X"a5",
X"54",
X"cd",
X"bf",
X"02",
X"90",
X"f4",
X"a2",
X"00",
X"f0",
X"ee",
X"c6",
X"55",
X"a5",
X"55",
X"30",
X"04",
X"c5",
X"52",
X"b0",
X"04",
X"a5",
X"53",
X"85",
X"55",
X"4c",
X"8e",
X"f8",
X"e6",
X"55",
X"a5",
X"55",
X"c5",
X"53",
X"90",
X"f5",
X"f0",
X"f3",
X"a5",
X"52",
X"4c",
X"0c",
X"f4",
X"20",
X"a6",
X"f9",
X"a4",
X"64",
X"a9",
X"00",
X"85",
X"64",
X"91",
X"64",
X"c8",
X"d0",
X"fb",
X"e6",
X"65",
X"a6",
X"65",
X"e4",
X"6a",
X"90",
X"f3",
X"a9",
X"ff",
X"99",
X"b2",
X"02",
X"c8",
X"c0",
X"04",
X"90",
X"f8",
X"20",
X"97",
X"f9",
X"85",
X"63",
X"85",
X"6d",
X"a9",
X"00",
X"85",
X"54",
X"85",
X"56",
X"85",
X"6c",
X"60",
X"a5",
X"63",
X"c5",
X"52",
X"f0",
X"21",
X"a5",
X"55",
X"c5",
X"52",
X"d0",
X"03",
X"20",
X"23",
X"f9",
X"20",
X"00",
X"f4",
X"a5",
X"55",
X"c5",
X"53",
X"d0",
X"07",
X"a5",
X"54",
X"f0",
X"03",
X"20",
X"e6",
X"f3",
X"a9",
X"20",
X"8d",
X"fb",
X"02",
X"20",
X"ca",
X"f1",
X"4c",
X"8e",
X"f8",
X"20",
X"11",
X"f4",
X"a5",
X"55",
X"c5",
X"52",
X"d0",
X"08",
X"20",
X"65",
X"f6",
X"20",
X"58",
X"f7",
X"b0",
X"07",
X"a5",
X"63",
X"20",
X"5d",
X"f7",
X"90",
X"e8",
X"4c",
X"8e",
X"f8",
X"a5",
X"63",
X"4c",
X"3e",
X"f7",
X"a5",
X"63",
X"4c",
X"4a",
X"f7",
X"20",
X"4c",
X"f9",
X"20",
X"8f",
X"f1",
X"85",
X"7d",
X"a9",
X"00",
X"8d",
X"bb",
X"02",
X"20",
X"e9",
X"f1",
X"a5",
X"63",
X"48",
X"20",
X"12",
X"f6",
X"68",
X"c5",
X"63",
X"b0",
X"0c",
X"a5",
X"7d",
X"48",
X"20",
X"8f",
X"f1",
X"85",
X"7d",
X"68",
X"4c",
X"ac",
X"f4",
X"20",
X"57",
X"f9",
X"ce",
X"bb",
X"02",
X"30",
X"04",
X"c6",
X"54",
X"d0",
X"f7",
X"4c",
X"8e",
X"f8",
X"20",
X"4c",
X"f9",
X"20",
X"ac",
X"f5",
X"a5",
X"64",
X"85",
X"68",
X"a5",
X"65",
X"85",
X"69",
X"a5",
X"63",
X"48",
X"20",
X"0a",
X"f6",
X"68",
X"c5",
X"63",
X"b0",
X"10",
X"a5",
X"54",
X"cd",
X"bf",
X"02",
X"b0",
X"09",
X"20",
X"8f",
X"f1",
X"a0",
X"00",
X"91",
X"68",
X"f0",
X"da",
X"a0",
X"00",
X"98",
X"91",
X"68",
X"20",
X"18",
X"f9",
X"20",
X"57",
X"f9",
X"4c",
X"8e",
X"f8",
X"38",
X"20",
X"c2",
X"f7",
X"a5",
X"52",
X"85",
X"55",
X"20",
X"ac",
X"f5",
X"20",
X"8e",
X"f7",
X"20",
X"e2",
X"f7",
X"4c",
X"8e",
X"f8",
X"20",
X"8e",
X"f8",
X"a4",
X"51",
X"84",
X"54",
X"a4",
X"54",
X"98",
X"38",
X"20",
X"5b",
X"f7",
X"08",
X"98",
X"18",
X"69",
X"78",
X"28",
X"20",
X"3c",
X"f7",
X"c8",
X"c0",
X"18",
X"d0",
X"ed",
X"ad",
X"b4",
X"02",
X"09",
X"01",
X"8d",
X"b4",
X"02",
X"a9",
X"00",
X"85",
X"55",
X"20",
X"ac",
X"f5",
X"20",
X"2a",
X"f8",
X"20",
X"58",
X"f7",
X"90",
X"d4",
X"4c",
X"1b",
X"f4",
X"a0",
X"20",
X"20",
X"83",
X"f9",
X"88",
X"10",
X"fa",
X"60",
X"20",
X"40",
X"f4",
X"4c",
X"e6",
X"f3",
X"a9",
X"02",
X"d0",
X"11",
X"ac",
X"6e",
X"02",
X"f0",
X"02",
X"09",
X"20",
X"a4",
X"4c",
X"30",
X"2b",
X"a0",
X"00",
X"91",
X"64",
X"a9",
X"01",
X"8d",
X"9e",
X"02",
X"a5",
X"4c",
X"30",
X"1e",
X"a5",
X"64",
X"38",
X"ed",
X"9e",
X"02",
X"85",
X"64",
X"b0",
X"02",
X"c6",
X"65",
X"a5",
X"0f",
X"c5",
X"65",
X"90",
X"0c",
X"d0",
X"06",
X"a5",
X"0e",
X"c5",
X"64",
X"90",
X"04",
X"a9",
X"93",
X"85",
X"4c",
X"60",
X"a9",
X"02",
X"20",
X"70",
X"f5",
X"a9",
X"a2",
X"20",
X"70",
X"f5",
X"ca",
X"60",
X"a2",
X"01",
X"86",
X"66",
X"ca",
X"86",
X"65",
X"a5",
X"54",
X"0a",
X"26",
X"65",
X"0a",
X"26",
X"65",
X"65",
X"54",
X"85",
X"64",
X"90",
X"02",
X"e6",
X"65",
X"a4",
X"57",
X"be",
X"6d",
X"ee",
X"06",
X"64",
X"26",
X"65",
X"ca",
X"d0",
X"f9",
X"a5",
X"56",
X"4a",
X"a5",
X"55",
X"be",
X"9d",
X"ee",
X"f0",
X"06",
X"6a",
X"06",
X"66",
X"ca",
X"d0",
X"fa",
X"65",
X"64",
X"90",
X"02",
X"e6",
X"65",
X"18",
X"65",
X"58",
X"85",
X"64",
X"85",
X"5e",
X"a5",
X"65",
X"65",
X"59",
X"85",
X"65",
X"85",
X"5f",
X"be",
X"9d",
X"ee",
X"bd",
X"04",
X"fb",
X"25",
X"55",
X"65",
X"66",
X"a8",
X"b9",
X"ac",
X"ee",
X"8d",
X"a0",
X"02",
X"85",
X"6f",
X"a0",
X"00",
X"60",
X"a9",
X"00",
X"f0",
X"02",
X"a9",
X"9b",
X"85",
X"7d",
X"e6",
X"63",
X"e6",
X"55",
X"d0",
X"02",
X"e6",
X"56",
X"a5",
X"55",
X"a6",
X"57",
X"dd",
X"7d",
X"ee",
X"f0",
X"0a",
X"e0",
X"00",
X"d0",
X"e2",
X"c5",
X"53",
X"f0",
X"de",
X"90",
X"dc",
X"e0",
X"08",
X"d0",
X"04",
X"a5",
X"56",
X"f0",
X"d4",
X"a5",
X"57",
X"d0",
X"2c",
X"a5",
X"63",
X"c9",
X"51",
X"90",
X"0a",
X"a5",
X"7d",
X"f0",
X"22",
X"20",
X"61",
X"f6",
X"4c",
X"ab",
X"f6",
X"20",
X"65",
X"f6",
X"a5",
X"54",
X"18",
X"69",
X"78",
X"20",
X"5d",
X"f7",
X"90",
X"08",
X"a5",
X"7d",
X"f0",
X"04",
X"18",
X"20",
X"0d",
X"f5",
X"4c",
X"8e",
X"f8",
X"a9",
X"9b",
X"85",
X"7d",
X"20",
X"97",
X"f9",
X"a9",
X"00",
X"85",
X"56",
X"e6",
X"54",
X"a6",
X"57",
X"a0",
X"18",
X"24",
X"7b",
X"10",
X"05",
X"a0",
X"04",
X"98",
X"d0",
X"03",
X"bd",
X"8d",
X"ee",
X"c5",
X"54",
X"d0",
X"29",
X"8c",
X"9d",
X"02",
X"8a",
X"d0",
X"23",
X"a5",
X"7d",
X"f0",
X"1f",
X"c9",
X"9b",
X"f0",
X"01",
X"18",
X"20",
X"f7",
X"f7",
X"ee",
X"bb",
X"02",
X"c6",
X"6c",
X"10",
X"02",
X"e6",
X"6c",
X"ce",
X"9d",
X"02",
X"ad",
X"b2",
X"02",
X"38",
X"10",
X"eb",
X"ad",
X"9d",
X"02",
X"85",
X"54",
X"4c",
X"8e",
X"f8",
X"38",
X"b5",
X"70",
X"e5",
X"74",
X"95",
X"70",
X"b5",
X"71",
X"e5",
X"75",
X"95",
X"71",
X"60",
X"ad",
X"bf",
X"02",
X"c9",
X"04",
X"f0",
X"07",
X"a5",
X"57",
X"f0",
X"03",
X"20",
X"94",
X"ef",
X"a9",
X"27",
X"c5",
X"53",
X"b0",
X"02",
X"85",
X"53",
X"a6",
X"57",
X"bd",
X"8d",
X"ee",
X"c5",
X"54",
X"90",
X"2a",
X"f0",
X"28",
X"e0",
X"08",
X"d0",
X"0a",
X"a5",
X"56",
X"f0",
X"13",
X"c9",
X"01",
X"d0",
X"1c",
X"f0",
X"04",
X"a5",
X"56",
X"d0",
X"16",
X"bd",
X"7d",
X"ee",
X"c5",
X"55",
X"90",
X"0f",
X"f0",
X"0d",
X"a9",
X"01",
X"85",
X"4c",
X"a9",
X"80",
X"a6",
X"11",
X"85",
X"11",
X"f0",
X"06",
X"60",
X"20",
X"40",
X"f4",
X"a9",
X"8d",
X"85",
X"4c",
X"68",
X"68",
X"a5",
X"7b",
X"10",
X"03",
X"4c",
X"62",
X"f9",
X"4c",
X"1e",
X"f2",
X"a0",
X"00",
X"a5",
X"5f",
X"f0",
X"04",
X"a5",
X"5d",
X"91",
X"5e",
X"60",
X"48",
X"29",
X"07",
X"aa",
X"bd",
X"b4",
X"ee",
X"85",
X"6e",
X"68",
X"4a",
X"4a",
X"4a",
X"aa",
X"60",
X"2e",
X"b4",
X"02",
X"2e",
X"b3",
X"02",
X"2e",
X"b2",
X"02",
X"60",
X"90",
X"0c",
X"20",
X"23",
X"f7",
X"bd",
X"a3",
X"02",
X"05",
X"6e",
X"9d",
X"a3",
X"02",
X"60",
X"20",
X"23",
X"f7",
X"a5",
X"6e",
X"49",
X"ff",
X"3d",
X"a3",
X"02",
X"9d",
X"a3",
X"02",
X"60",
X"a5",
X"54",
X"18",
X"69",
X"78",
X"20",
X"23",
X"f7",
X"18",
X"bd",
X"a3",
X"02",
X"25",
X"6e",
X"f0",
X"01",
X"38",
X"60",
X"ad",
X"fa",
X"02",
X"a4",
X"57",
X"c0",
X"0e",
X"b0",
X"17",
X"c0",
X"0c",
X"b0",
X"04",
X"c0",
X"03",
X"b0",
X"0f",
X"2a",
X"2a",
X"2a",
X"2a",
X"29",
X"03",
X"aa",
X"ad",
X"fa",
X"02",
X"29",
X"9f",
X"1d",
X"4d",
X"fb",
X"8d",
X"fb",
X"02",
X"60",
X"a6",
X"6a",
X"ca",
X"86",
X"69",
X"86",
X"67",
X"a9",
X"b0",
X"85",
X"68",
X"a9",
X"d8",
X"85",
X"66",
X"a6",
X"54",
X"e8",
X"ec",
X"bf",
X"02",
X"f0",
X"e8",
X"a0",
X"27",
X"b1",
X"68",
X"91",
X"66",
X"88",
X"10",
X"f9",
X"38",
X"a5",
X"68",
X"85",
X"66",
X"e9",
X"28",
X"85",
X"68",
X"a5",
X"69",
X"85",
X"67",
X"e9",
X"00",
X"85",
X"69",
X"4c",
X"9f",
X"f7",
X"08",
X"a0",
X"16",
X"98",
X"20",
X"5a",
X"f7",
X"08",
X"98",
X"18",
X"69",
X"79",
X"28",
X"20",
X"3c",
X"f7",
X"88",
X"30",
X"04",
X"c4",
X"54",
X"b0",
X"ec",
X"a5",
X"54",
X"18",
X"69",
X"78",
X"28",
X"4c",
X"3c",
X"f7",
X"a5",
X"52",
X"85",
X"55",
X"20",
X"ac",
X"f5",
X"38",
X"a5",
X"53",
X"e5",
X"52",
X"a8",
X"a9",
X"00",
X"91",
X"64",
X"88",
X"10",
X"fb",
X"60",
X"20",
X"32",
X"f7",
X"ad",
X"6e",
X"02",
X"f0",
X"28",
X"ad",
X"6c",
X"02",
X"d0",
X"fb",
X"a9",
X"08",
X"8d",
X"6c",
X"02",
X"ad",
X"6c",
X"02",
X"c9",
X"01",
X"d0",
X"f9",
X"ad",
X"0b",
X"d4",
X"c9",
X"40",
X"b0",
X"f9",
X"a2",
X"0d",
X"ad",
X"bf",
X"02",
X"c9",
X"04",
X"d0",
X"02",
X"a2",
X"70",
X"ec",
X"0b",
X"d4",
X"b0",
X"fb",
X"20",
X"a6",
X"f9",
X"a5",
X"64",
X"a6",
X"65",
X"e8",
X"e4",
X"6a",
X"f0",
X"06",
X"38",
X"e9",
X"10",
X"4c",
X"2e",
X"f8",
X"69",
X"27",
X"d0",
X"0a",
X"a6",
X"65",
X"e8",
X"e4",
X"6a",
X"f0",
X"38",
X"18",
X"69",
X"10",
X"a8",
X"85",
X"7e",
X"38",
X"a5",
X"64",
X"e5",
X"7e",
X"85",
X"64",
X"b0",
X"02",
X"c6",
X"65",
X"a5",
X"64",
X"18",
X"69",
X"28",
X"85",
X"7e",
X"a5",
X"65",
X"69",
X"00",
X"85",
X"7f",
X"b1",
X"7e",
X"91",
X"64",
X"c8",
X"d0",
X"f9",
X"a0",
X"10",
X"a5",
X"64",
X"c9",
X"d8",
X"f0",
X"0b",
X"18",
X"69",
X"f0",
X"85",
X"64",
X"90",
X"dd",
X"e6",
X"65",
X"d0",
X"d9",
X"a6",
X"6a",
X"ca",
X"86",
X"7f",
X"a2",
X"d8",
X"86",
X"7e",
X"a9",
X"00",
X"a0",
X"27",
X"91",
X"7e",
X"88",
X"10",
X"fb",
X"a9",
X"00",
X"85",
X"63",
X"a5",
X"54",
X"85",
X"51",
X"a5",
X"51",
X"20",
X"5a",
X"f7",
X"b0",
X"0c",
X"a5",
X"63",
X"18",
X"69",
X"28",
X"85",
X"63",
X"c6",
X"51",
X"4c",
X"96",
X"f8",
X"18",
X"a5",
X"63",
X"65",
X"55",
X"85",
X"63",
X"60",
X"20",
X"4c",
X"f9",
X"a5",
X"63",
X"48",
X"a5",
X"6c",
X"85",
X"54",
X"a5",
X"6d",
X"85",
X"55",
X"a9",
X"01",
X"85",
X"6b",
X"a2",
X"17",
X"a5",
X"7b",
X"10",
X"02",
X"a2",
X"03",
X"e4",
X"54",
X"d0",
X"0b",
X"a5",
X"55",
X"c5",
X"53",
X"d0",
X"05",
X"e6",
X"6b",
X"4c",
X"ea",
X"f8",
X"20",
X"0a",
X"f6",
X"e6",
X"6b",
X"a5",
X"63",
X"c5",
X"52",
X"d0",
X"de",
X"c6",
X"54",
X"20",
X"00",
X"f4",
X"20",
X"8f",
X"f1",
X"d0",
X"17",
X"c6",
X"6b",
X"a5",
X"63",
X"c5",
X"52",
X"f0",
X"0f",
X"20",
X"00",
X"f4",
X"a5",
X"55",
X"c5",
X"53",
X"d0",
X"02",
X"c6",
X"54",
X"a5",
X"6b",
X"d0",
X"e4",
X"68",
X"85",
X"63",
X"4c",
X"57",
X"f9",
X"20",
X"8e",
X"f8",
X"a5",
X"51",
X"85",
X"6c",
X"a5",
X"52",
X"85",
X"6d",
X"60",
X"a5",
X"63",
X"c5",
X"52",
X"d0",
X"02",
X"c6",
X"54",
X"20",
X"8e",
X"f8",
X"a5",
X"63",
X"c5",
X"52",
X"f0",
X"ee",
X"20",
X"ac",
X"f5",
X"a5",
X"53",
X"38",
X"e5",
X"52",
X"a8",
X"b1",
X"64",
X"d0",
X"e1",
X"88",
X"10",
X"f9",
X"4c",
X"27",
X"f5",
X"a2",
X"2d",
X"bd",
X"0d",
X"fb",
X"cd",
X"fb",
X"02",
X"f0",
X"05",
X"ca",
X"ca",
X"ca",
X"10",
X"f3",
X"60",
X"a2",
X"02",
X"b5",
X"54",
X"9d",
X"b8",
X"02",
X"ca",
X"10",
X"f8",
X"60",
X"a2",
X"02",
X"bd",
X"b8",
X"02",
X"95",
X"54",
X"ca",
X"10",
X"f8",
X"60",
X"ad",
X"bf",
X"02",
X"c9",
X"18",
X"f0",
X"17",
X"a2",
X"0b",
X"b5",
X"54",
X"48",
X"bd",
X"90",
X"02",
X"95",
X"54",
X"68",
X"9d",
X"90",
X"02",
X"ca",
X"10",
X"f1",
X"a5",
X"7b",
X"49",
X"ff",
X"85",
X"7b",
X"4c",
X"1e",
X"f2",
X"a2",
X"7e",
X"48",
X"8e",
X"1f",
X"d0",
X"ad",
X"0b",
X"d4",
X"cd",
X"0b",
X"d4",
X"f0",
X"fb",
X"ca",
X"ca",
X"10",
X"f1",
X"68",
X"60",
X"a9",
X"00",
X"a6",
X"7b",
X"d0",
X"04",
X"a6",
X"57",
X"d0",
X"02",
X"a5",
X"52",
X"85",
X"55",
X"60",
X"a5",
X"58",
X"85",
X"64",
X"a5",
X"59",
X"85",
X"65",
X"60",
X"a2",
X"00",
X"a5",
X"22",
X"c9",
X"11",
X"f0",
X"08",
X"c9",
X"12",
X"f0",
X"03",
X"a0",
X"84",
X"60",
X"e8",
X"8e",
X"b7",
X"02",
X"a5",
X"54",
X"8d",
X"f5",
X"02",
X"a5",
X"55",
X"8d",
X"f6",
X"02",
X"a5",
X"56",
X"8d",
X"f7",
X"02",
X"a9",
X"01",
X"8d",
X"f8",
X"02",
X"8d",
X"f9",
X"02",
X"38",
X"ad",
X"f5",
X"02",
X"e5",
X"5a",
X"85",
X"76",
X"b0",
X"0e",
X"a9",
X"ff",
X"8d",
X"f8",
X"02",
X"a5",
X"76",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"85",
X"76",
X"38",
X"ad",
X"f6",
X"02",
X"e5",
X"5b",
X"85",
X"77",
X"ad",
X"f7",
X"02",
X"e5",
X"5c",
X"85",
X"78",
X"b0",
X"17",
X"a9",
X"ff",
X"8d",
X"f9",
X"02",
X"a5",
X"77",
X"49",
X"ff",
X"85",
X"77",
X"a5",
X"78",
X"49",
X"ff",
X"85",
X"78",
X"e6",
X"77",
X"d0",
X"02",
X"e6",
X"78",
X"a2",
X"02",
X"a0",
X"00",
X"84",
X"73",
X"98",
X"95",
X"70",
X"b5",
X"5a",
X"95",
X"54",
X"ca",
X"10",
X"f6",
X"a5",
X"77",
X"e8",
X"a8",
X"a5",
X"78",
X"85",
X"7f",
X"85",
X"75",
X"d0",
X"0b",
X"a5",
X"77",
X"c5",
X"76",
X"b0",
X"05",
X"a5",
X"76",
X"a2",
X"02",
X"a8",
X"98",
X"85",
X"7e",
X"85",
X"74",
X"48",
X"a5",
X"75",
X"4a",
X"68",
X"6a",
X"95",
X"70",
X"a5",
X"7e",
X"05",
X"7f",
X"d0",
X"03",
X"4c",
X"01",
X"fb",
X"18",
X"a5",
X"70",
X"65",
X"76",
X"85",
X"70",
X"90",
X"02",
X"e6",
X"71",
X"a5",
X"71",
X"c5",
X"75",
X"90",
X"15",
X"d0",
X"06",
X"a5",
X"70",
X"c5",
X"74",
X"90",
X"0d",
X"18",
X"a5",
X"54",
X"6d",
X"f8",
X"02",
X"85",
X"54",
X"a2",
X"00",
X"20",
X"ae",
X"f6",
X"18",
X"a5",
X"72",
X"65",
X"77",
X"85",
X"72",
X"a5",
X"73",
X"65",
X"78",
X"85",
X"73",
X"c5",
X"75",
X"90",
X"28",
X"d0",
X"06",
X"a5",
X"72",
X"c5",
X"74",
X"90",
X"20",
X"2c",
X"f9",
X"02",
X"10",
X"10",
X"c6",
X"55",
X"a5",
X"55",
X"c9",
X"ff",
X"d0",
X"0e",
X"a5",
X"56",
X"f0",
X"0a",
X"c6",
X"56",
X"10",
X"06",
X"e6",
X"55",
X"d0",
X"02",
X"e6",
X"56",
X"a2",
X"02",
X"20",
X"ae",
X"f6",
X"20",
X"ca",
X"f6",
X"20",
X"ca",
X"f1",
X"ad",
X"b7",
X"02",
X"f0",
X"2f",
X"20",
X"4c",
X"f9",
X"ad",
X"fb",
X"02",
X"8d",
X"bc",
X"02",
X"a5",
X"54",
X"48",
X"20",
X"12",
X"f6",
X"68",
X"85",
X"54",
X"20",
X"ca",
X"f6",
X"20",
X"8f",
X"f1",
X"d0",
X"0c",
X"ad",
X"fd",
X"02",
X"8d",
X"fb",
X"02",
X"20",
X"ca",
X"f1",
X"4c",
X"c9",
X"fa",
X"ad",
X"bc",
X"02",
X"8d",
X"fb",
X"02",
X"20",
X"57",
X"f9",
X"38",
X"a5",
X"7e",
X"e9",
X"01",
X"85",
X"7e",
X"a5",
X"7f",
X"e9",
X"00",
X"85",
X"7f",
X"30",
X"03",
X"4c",
X"4d",
X"fa",
X"4c",
X"1e",
X"f2",
X"00",
X"01",
X"03",
X"07",
X"28",
X"ca",
X"94",
X"46",
X"00",
X"1b",
X"e0",
X"f3",
X"1c",
X"e6",
X"f3",
X"1d",
X"f3",
X"f3",
X"1e",
X"00",
X"f4",
X"1f",
X"11",
X"f4",
X"7d",
X"20",
X"f4",
X"7e",
X"50",
X"f4",
X"7f",
X"7a",
X"f4",
X"9b",
X"61",
X"f6",
X"9c",
X"20",
X"f5",
X"9d",
X"0c",
X"f5",
X"9e",
X"9a",
X"f4",
X"9f",
X"95",
X"f4",
X"fd",
X"56",
X"f5",
X"fe",
X"d5",
X"f4",
X"ff",
X"9f",
X"f4",
X"1c",
X"40",
X"f4",
X"1d",
X"5f",
X"f5",
X"1e",
X"1b",
X"f4",
X"1f",
X"0a",
X"f4",
X"40",
X"00",
X"20",
X"60",
X"20",
X"40",
X"00",
X"60",
X"6c",
X"6a",
X"3b",
X"8a",
X"8b",
X"6b",
X"2b",
X"2a",
X"6f",
X"80",
X"70",
X"75",
X"9b",
X"69",
X"2d",
X"3d",
X"76",
X"80",
X"63",
X"8c",
X"8d",
X"62",
X"78",
X"7a",
X"34",
X"80",
X"33",
X"36",
X"1b",
X"35",
X"32",
X"31",
X"2c",
X"20",
X"2e",
X"6e",
X"80",
X"6d",
X"2f",
X"81",
X"72",
X"80",
X"65",
X"79",
X"7f",
X"74",
X"77",
X"71",
X"39",
X"80",
X"30",
X"37",
X"7e",
X"38",
X"3c",
X"3e",
X"66",
X"68",
X"64",
X"80",
X"82",
X"67",
X"73",
X"61",
X"4c",
X"4a",
X"3a",
X"8a",
X"8b",
X"4b",
X"5c",
X"5e",
X"4f",
X"80",
X"50",
X"55",
X"9b",
X"49",
X"5f",
X"7c",
X"56",
X"80",
X"43",
X"8c",
X"8d",
X"42",
X"58",
X"5a",
X"24",
X"80",
X"23",
X"26",
X"1b",
X"25",
X"22",
X"21",
X"5b",
X"20",
X"5d",
X"4e",
X"80",
X"4d",
X"3f",
X"81",
X"52",
X"80",
X"45",
X"59",
X"9f",
X"54",
X"57",
X"51",
X"28",
X"80",
X"29",
X"27",
X"9c",
X"40",
X"7d",
X"9d",
X"46",
X"48",
X"44",
X"80",
X"83",
X"47",
X"53",
X"41",
X"0c",
X"0a",
X"7b",
X"80",
X"80",
X"0b",
X"1e",
X"1f",
X"0f",
X"80",
X"10",
X"15",
X"9b",
X"09",
X"1c",
X"1d",
X"16",
X"80",
X"03",
X"89",
X"80",
X"02",
X"18",
X"1a",
X"80",
X"80",
X"85",
X"80",
X"1b",
X"80",
X"fd",
X"80",
X"00",
X"20",
X"60",
X"0e",
X"80",
X"0d",
X"80",
X"81",
X"12",
X"80",
X"05",
X"19",
X"9e",
X"14",
X"17",
X"11",
X"80",
X"80",
X"80",
X"80",
X"fe",
X"80",
X"7d",
X"ff",
X"06",
X"08",
X"04",
X"80",
X"84",
X"07",
X"13",
X"01",
X"1c",
X"1d",
X"1e",
X"1f",
X"8e",
X"8f",
X"90",
X"91",
X"8a",
X"48",
X"98",
X"48",
X"ac",
X"01",
X"d3",
X"ad",
X"09",
X"d2",
X"cd",
X"f2",
X"02",
X"d0",
X"05",
X"ae",
X"f1",
X"02",
X"d0",
X"49",
X"ae",
X"6d",
X"02",
X"c9",
X"83",
X"d0",
X"13",
X"8a",
X"49",
X"ff",
X"8d",
X"6d",
X"02",
X"d0",
X"05",
X"98",
X"09",
X"04",
X"d0",
X"03",
X"98",
X"29",
X"fb",
X"a8",
X"b0",
X"26",
X"8a",
X"d0",
X"3d",
X"ad",
X"09",
X"d2",
X"aa",
X"c9",
X"9f",
X"d0",
X"0a",
X"ad",
X"ff",
X"02",
X"49",
X"ff",
X"8d",
X"ff",
X"02",
X"b0",
X"11",
X"29",
X"3f",
X"c9",
X"11",
X"d0",
X"2e",
X"8e",
X"dc",
X"02",
X"f0",
X"06",
X"8e",
X"fc",
X"02",
X"8e",
X"f2",
X"02",
X"a9",
X"03",
X"8d",
X"f1",
X"02",
X"a9",
X"00",
X"85",
X"4d",
X"ad",
X"d9",
X"02",
X"8d",
X"2b",
X"02",
X"ad",
X"2f",
X"02",
X"d0",
X"06",
X"ad",
X"dd",
X"02",
X"8d",
X"2f",
X"02",
X"8c",
X"01",
X"d3",
X"68",
X"a8",
X"68",
X"aa",
X"68",
X"40",
X"e0",
X"84",
X"f0",
X"21",
X"e0",
X"94",
X"d0",
X"cf",
X"ad",
X"f4",
X"02",
X"ae",
X"6b",
X"02",
X"8d",
X"6b",
X"02",
X"8e",
X"f4",
X"02",
X"e0",
X"cc",
X"f0",
X"06",
X"98",
X"09",
X"08",
X"a8",
X"d0",
X"bf",
X"98",
X"29",
X"f7",
X"a8",
X"4c",
X"6d",
X"fc",
X"ad",
X"2f",
X"02",
X"f0",
X"cd",
X"8d",
X"dd",
X"02",
X"a9",
X"00",
X"8d",
X"2f",
X"02",
X"f0",
X"c3",
X"48",
X"ad",
X"c6",
X"02",
X"4d",
X"4f",
X"00",
X"2d",
X"4e",
X"00",
X"8d",
X"0a",
X"d4",
X"8d",
X"17",
X"d0",
X"68",
X"40",
X"00",
X"00",
X"4c",
X"83",
X"f9",
X"a9",
X"cc",
X"8d",
X"ee",
X"02",
X"a9",
X"05",
X"8d",
X"ef",
X"02",
X"60",
X"a5",
X"2b",
X"85",
X"3e",
X"a5",
X"2a",
X"29",
X"0c",
X"c9",
X"04",
X"f0",
X"05",
X"c9",
X"08",
X"f0",
X"3e",
X"60",
X"a9",
X"00",
X"8d",
X"89",
X"02",
X"85",
X"3f",
X"a9",
X"01",
X"20",
X"fc",
X"fd",
X"30",
X"29",
X"a9",
X"34",
X"8d",
X"02",
X"d3",
X"a6",
X"62",
X"bc",
X"93",
X"fe",
X"bd",
X"91",
X"fe",
X"aa",
X"a9",
X"03",
X"8d",
X"2a",
X"02",
X"20",
X"5c",
X"e4",
X"ad",
X"2a",
X"02",
X"d0",
X"fb",
X"a9",
X"80",
X"85",
X"3d",
X"8d",
X"8a",
X"02",
X"4c",
X"77",
X"fd",
X"a0",
X"80",
X"c6",
X"11",
X"a9",
X"00",
X"8d",
X"89",
X"02",
X"60",
X"a9",
X"80",
X"8d",
X"89",
X"02",
X"a9",
X"02",
X"20",
X"fc",
X"fd",
X"30",
X"ee",
X"a9",
X"cc",
X"8d",
X"04",
X"d2",
X"a9",
X"05",
X"8d",
X"06",
X"d2",
X"a9",
X"60",
X"8d",
X"00",
X"03",
X"20",
X"68",
X"e4",
X"a9",
X"34",
X"8d",
X"02",
X"d3",
X"a6",
X"62",
X"bc",
X"8f",
X"fe",
X"bd",
X"8d",
X"fe",
X"aa",
X"a9",
X"03",
X"20",
X"5c",
X"e4",
X"a9",
X"ff",
X"8d",
X"2a",
X"02",
X"a5",
X"11",
X"f0",
X"bc",
X"ad",
X"2a",
X"02",
X"d0",
X"f7",
X"a9",
X"00",
X"85",
X"3d",
X"a0",
X"01",
X"60",
X"a5",
X"3f",
X"30",
X"33",
X"a6",
X"3d",
X"ec",
X"8a",
X"02",
X"f0",
X"08",
X"bd",
X"00",
X"04",
X"e6",
X"3d",
X"a0",
X"01",
X"60",
X"a9",
X"52",
X"20",
X"3f",
X"fe",
X"98",
X"30",
X"f7",
X"a9",
X"00",
X"85",
X"3d",
X"a2",
X"80",
X"ad",
X"ff",
X"03",
X"c9",
X"fe",
X"f0",
X"0d",
X"c9",
X"fa",
X"d0",
X"03",
X"ae",
X"7f",
X"04",
X"8e",
X"8a",
X"02",
X"4c",
X"7a",
X"fd",
X"c6",
X"3f",
X"a0",
X"88",
X"60",
X"a6",
X"3d",
X"9d",
X"00",
X"04",
X"e6",
X"3d",
X"a0",
X"01",
X"e0",
X"7f",
X"f0",
X"01",
X"60",
X"a9",
X"fc",
X"20",
X"7c",
X"fe",
X"a9",
X"00",
X"85",
X"3d",
X"60",
X"a0",
X"01",
X"60",
X"ad",
X"89",
X"02",
X"30",
X"08",
X"a0",
X"01",
X"a9",
X"3c",
X"8d",
X"02",
X"d3",
X"60",
X"a6",
X"3d",
X"f0",
X"0a",
X"8e",
X"7f",
X"04",
X"a9",
X"fa",
X"20",
X"7c",
X"fe",
X"30",
X"ec",
X"a2",
X"7f",
X"a9",
X"00",
X"9d",
X"00",
X"04",
X"ca",
X"10",
X"fa",
X"a9",
X"fe",
X"20",
X"7c",
X"fe",
X"4c",
X"d6",
X"fd",
X"85",
X"40",
X"a5",
X"14",
X"18",
X"a6",
X"62",
X"7d",
X"95",
X"fe",
X"aa",
X"a9",
X"ff",
X"8d",
X"1f",
X"d0",
X"a9",
X"00",
X"a0",
X"f0",
X"88",
X"d0",
X"fd",
X"8d",
X"1f",
X"d0",
X"a0",
X"f0",
X"88",
X"d0",
X"fd",
X"e4",
X"14",
X"d0",
X"e8",
X"c6",
X"40",
X"f0",
X"0e",
X"8a",
X"18",
X"a6",
X"62",
X"7d",
X"97",
X"fe",
X"aa",
X"e4",
X"14",
X"d0",
X"fc",
X"f0",
X"cd",
X"20",
X"36",
X"fe",
X"98",
X"60",
X"ad",
X"25",
X"e4",
X"48",
X"ad",
X"24",
X"e4",
X"48",
X"60",
X"8d",
X"02",
X"03",
X"a9",
X"00",
X"8d",
X"09",
X"03",
X"a9",
X"83",
X"8d",
X"08",
X"03",
X"a9",
X"03",
X"8d",
X"05",
X"03",
X"a9",
X"fd",
X"8d",
X"04",
X"03",
X"a9",
X"60",
X"8d",
X"00",
X"03",
X"a9",
X"00",
X"8d",
X"01",
X"03",
X"a9",
X"23",
X"8d",
X"06",
X"03",
X"ad",
X"02",
X"03",
X"a0",
X"40",
X"c9",
X"52",
X"f0",
X"02",
X"a0",
X"80",
X"8c",
X"03",
X"03",
X"a5",
X"3e",
X"8d",
X"0b",
X"03",
X"20",
X"59",
X"e4",
X"60",
X"8d",
X"ff",
X"03",
X"a9",
X"55",
X"8d",
X"fd",
X"03",
X"8d",
X"fe",
X"03",
X"a9",
X"57",
X"20",
X"3f",
X"fe",
X"60",
X"04",
X"03",
X"80",
X"c0",
X"02",
X"01",
X"40",
X"e0",
X"1e",
X"19",
X"0a",
X"08",
X"a9",
X"1e",
X"8d",
X"14",
X"03",
X"60",
X"ea",
X"02",
X"c0",
X"03",
X"a9",
X"04",
X"8d",
X"df",
X"02",
X"ae",
X"9f",
X"fe",
X"ac",
X"a0",
X"fe",
X"a9",
X"53",
X"8d",
X"02",
X"03",
X"8d",
X"0a",
X"03",
X"20",
X"14",
X"ff",
X"20",
X"59",
X"e4",
X"30",
X"03",
X"20",
X"44",
X"ff",
X"60",
X"20",
X"a3",
X"fe",
X"a9",
X"00",
X"8d",
X"de",
X"02",
X"60",
X"48",
X"bd",
X"41",
X"03",
X"85",
X"21",
X"20",
X"4b",
X"ff",
X"ae",
X"de",
X"02",
X"68",
X"9d",
X"c0",
X"03",
X"e8",
X"ec",
X"df",
X"02",
X"f0",
X"15",
X"8e",
X"de",
X"02",
X"c9",
X"9b",
X"f0",
X"03",
X"a0",
X"01",
X"60",
X"a9",
X"20",
X"9d",
X"c0",
X"03",
X"e8",
X"ec",
X"df",
X"02",
X"d0",
X"f7",
X"a9",
X"00",
X"8d",
X"de",
X"02",
X"ae",
X"a1",
X"fe",
X"ac",
X"a2",
X"fe",
X"20",
X"14",
X"ff",
X"4c",
X"59",
X"e4",
X"20",
X"4b",
X"ff",
X"a9",
X"9b",
X"ae",
X"de",
X"02",
X"d0",
X"dc",
X"a0",
X"01",
X"60",
X"8e",
X"04",
X"03",
X"8c",
X"05",
X"03",
X"a9",
X"40",
X"8d",
X"00",
X"03",
X"a5",
X"21",
X"8d",
X"01",
X"03",
X"a9",
X"80",
X"ae",
X"02",
X"03",
X"e0",
X"53",
X"d0",
X"02",
X"a9",
X"40",
X"8d",
X"03",
X"03",
X"ad",
X"df",
X"02",
X"8d",
X"08",
X"03",
X"a9",
X"00",
X"8d",
X"09",
X"03",
X"ad",
X"14",
X"03",
X"8d",
X"06",
X"03",
X"60",
X"ad",
X"ec",
X"02",
X"8d",
X"14",
X"03",
X"60",
X"a0",
X"57",
X"a5",
X"2b",
X"c9",
X"4e",
X"d0",
X"04",
X"a2",
X"28",
X"d0",
X"0e",
X"c9",
X"44",
X"d0",
X"04",
X"a2",
X"14",
X"d0",
X"06",
X"c9",
X"53",
X"d0",
X"0c",
X"a2",
X"1d",
X"8e",
X"df",
X"02",
X"8c",
X"02",
X"03",
X"8d",
X"0a",
X"03",
X"60",
X"a9",
X"4e",
X"d0",
X"dc",
X"a2",
X"00",
X"86",
X"8b",
X"86",
X"8c",
X"20",
X"a9",
X"ff",
X"e0",
X"0c",
X"d0",
X"f9",
X"ad",
X"00",
X"c0",
X"ae",
X"01",
X"c0",
X"c5",
X"8b",
X"d0",
X"06",
X"e4",
X"8c",
X"d0",
X"02",
X"18",
X"60",
X"38",
X"60",
X"a2",
X"00",
X"86",
X"8b",
X"86",
X"8c",
X"a2",
X"0c",
X"20",
X"a9",
X"ff",
X"20",
X"a9",
X"ff",
X"ad",
X"f8",
X"ff",
X"ae",
X"f9",
X"ff",
X"4c",
X"86",
X"ff",
X"a0",
X"00",
X"bd",
X"d7",
X"ff",
X"99",
X"9e",
X"00",
X"e8",
X"c8",
X"c0",
X"04",
X"d0",
X"f4",
X"a0",
X"00",
X"18",
X"b1",
X"9e",
X"65",
X"8b",
X"85",
X"8b",
X"90",
X"02",
X"e6",
X"8c",
X"e6",
X"9e",
X"d0",
X"02",
X"e6",
X"9f",
X"a5",
X"9e",
X"c5",
X"a0",
X"d0",
X"e9",
X"a5",
X"9f",
X"c5",
X"a1",
X"d0",
X"e3",
X"60",
X"02",
X"c0",
X"00",
X"d0",
X"00",
X"50",
X"00",
X"58",
X"00",
X"d8",
X"00",
X"e0",
X"00",
X"e0",
X"f8",
X"ff",
X"fa",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"10",
X"05",
X"83",
X"02",
X"42",
X"42",
X"00",
X"00",
X"01",
X"02",
X"8c",
X"6c",
X"18",
X"c0",
X"00",
X"c0",
X"2c",
X"c0"

);
        signal rdata:std_logic_vector(7 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
