-------------------------------------------------------------------------------
--
-- $Id: T80_MCode-c.vhd,v 1.1 2006/01/03 08:23:24 arnim Exp $
--
-------------------------------------------------------------------------------

configuration T80_MCode_rtl_c0 of T80_MCode is

  for rtl
  end for;

end T80_MCode_rtl_c0;
