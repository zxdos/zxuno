-------------------------------------------------------------------------------
--
-- FPGA Colecovision
--
-- $Id: cv_clock-c.vhd,v 1.2 2006/01/05 22:25:25 arnim Exp $
--
-------------------------------------------------------------------------------

configuration cv_clock_rtl_c0 of cv_clock is

  for rtl
  end for;

end cv_clock_rtl_c0;
