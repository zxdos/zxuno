-------------------------------------------------------------------------------
--
-- FPGA Colecovision
--
-- $Id: cv_ctrl-c.vhd,v 1.2 2006/01/05 22:25:25 arnim Exp $
--
-------------------------------------------------------------------------------

configuration cv_ctrl_rtl_c0 of cv_ctrl is

  for rtl
  end for;

end cv_ctrl_rtl_c0;
