-------------------------------------------------------------------------------
--
-- SNESpad controller core
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- $Id: snespad_ctrl-c.vhd,v 1.1 2004/10/05 17:01:27 arniml Exp $
--
-------------------------------------------------------------------------------

configuration snespad_ctrl_rtl_c0 of snespad_ctrl is

  for rtl
  end for;

end snespad_ctrl_rtl_c0;
