-- generated with romgen by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity VIC20_GAME_ROM is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of VIC20_GAME_ROM is


  type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"00",x"A0",x"09",x"A0",x"56",x"FF",x"41",x"30", -- 0x0000
    x"C3",x"C2",x"CD",x"78",x"20",x"8D",x"A6",x"A9", -- 0x0008
    x"00",x"85",x"EE",x"85",x"EB",x"85",x"EF",x"85", -- 0x0010
    x"EC",x"85",x"F0",x"85",x"ED",x"EA",x"EA",x"EA", -- 0x0018
    x"EA",x"AA",x"4C",x"46",x"AA",x"85",x"09",x"A9", -- 0x0020
    x"00",x"85",x"0A",x"06",x"09",x"26",x"0A",x"06", -- 0x0028
    x"09",x"26",x"0A",x"06",x"09",x"26",x"0A",x"A5", -- 0x0030
    x"0A",x"09",x"88",x"85",x"0A",x"4C",x"21",x"A7", -- 0x0038
    x"56",x"09",x"04",x"05",x"0F",x"0D",x"01",x"0E", -- 0x0040
    x"09",x"01",x"02",x"19",x"54",x"0F",x"0D",x"47", -- 0x0048
    x"12",x"09",x"0E",x"05",x"12",x"2C",x"34",x"3C", -- 0x0050
    x"44",x"4C",x"54",x"5C",x"64",x"6C",x"74",x"4C", -- 0x0058
    x"54",x"2C",x"34",x"3C",x"4C",x"54",x"5C",x"64", -- 0x0060
    x"6C",x"74",x"48",x"48",x"48",x"48",x"48",x"48", -- 0x0068
    x"48",x"48",x"48",x"48",x"50",x"50",x"58",x"58", -- 0x0070
    x"58",x"58",x"58",x"58",x"58",x"58",x"58",x"A5", -- 0x0078
    x"00",x"18",x"65",x"0D",x"85",x"00",x"A5",x"01", -- 0x0080
    x"69",x"00",x"85",x"01",x"60",x"20",x"0E",x"A1", -- 0x0088
    x"20",x"66",x"AD",x"20",x"77",x"AD",x"A9",x"00", -- 0x0090
    x"85",x"0D",x"85",x"0C",x"A9",x"FF",x"85",x"0F", -- 0x0098
    x"A2",x"14",x"20",x"A6",x"A8",x"95",x"B7",x"85", -- 0x00A0
    x"04",x"20",x"A6",x"A8",x"95",x"CC",x"85",x"05", -- 0x00A8
    x"BD",x"3E",x"A0",x"20",x"23",x"A0",x"CA",x"10", -- 0x00B0
    x"E9",x"A9",x"96",x"85",x"0C",x"A2",x"14",x"B5", -- 0x00B8
    x"B7",x"85",x"04",x"B5",x"CC",x"85",x"05",x"BD", -- 0x00C0
    x"3E",x"A0",x"20",x"23",x"A0",x"B5",x"B7",x"DD", -- 0x00C8
    x"53",x"A0",x"F0",x"09",x"90",x"05",x"D6",x"B7", -- 0x00D0
    x"4C",x"DB",x"A0",x"F6",x"B7",x"B5",x"CC",x"DD", -- 0x00D8
    x"68",x"A0",x"F0",x"09",x"90",x"05",x"D6",x"CC", -- 0x00E0
    x"4C",x"EB",x"A0",x"F6",x"CC",x"B5",x"B7",x"85", -- 0x00E8
    x"04",x"B5",x"CC",x"85",x"05",x"BD",x"3E",x"A0", -- 0x00F0
    x"20",x"23",x"A0",x"20",x"3B",x"A4",x"CA",x"10", -- 0x00F8
    x"BE",x"20",x"84",x"A8",x"29",x"20",x"F0",x"07", -- 0x0100
    x"C6",x"0C",x"D0",x"B1",x"4C",x"62",x"A1",x"60", -- 0x0108
    x"20",x"C0",x"AF",x"85",x"E7",x"20",x"07",x"A7", -- 0x0110
    x"A2",x"10",x"A9",x"00",x"95",x"48",x"CA",x"10", -- 0x0118
    x"F9",x"A2",x"07",x"A9",x"54",x"95",x"48",x"95", -- 0x0120
    x"59",x"8A",x"95",x"6A",x"CA",x"10",x"F4",x"A2", -- 0x0128
    x"50",x"8A",x"48",x"20",x"72",x"AB",x"E6",x"0C", -- 0x0130
    x"20",x"9A",x"A8",x"09",x"80",x"8D",x"0D",x"90", -- 0x0138
    x"68",x"AA",x"CA",x"D0",x"EC",x"20",x"C0",x"AF", -- 0x0140
    x"60",x"A6",x"EA",x"F0",x"FB",x"CA",x"A9",x"00", -- 0x0148
    x"85",x"04",x"A9",x"08",x"85",x"05",x"20",x"5A", -- 0x0150
    x"A9",x"A5",x"04",x"18",x"69",x"09",x"85",x"04", -- 0x0158
    x"CA",x"10",x"F3",x"60",x"A2",x"39",x"A9",x"00", -- 0x0160
    x"85",x"48",x"85",x"59",x"20",x"E0",x"A1",x"20", -- 0x0168
    x"E0",x"A1",x"A5",x"48",x"DD",x"F9",x"A1",x"F0", -- 0x0170
    x"09",x"B0",x"05",x"E6",x"48",x"4C",x"80",x"A1", -- 0x0178
    x"C6",x"48",x"A5",x"59",x"DD",x"33",x"A2",x"F0", -- 0x0180
    x"09",x"B0",x"05",x"E6",x"59",x"4C",x"90",x"A1", -- 0x0188
    x"C6",x"59",x"A5",x"48",x"DD",x"F9",x"A1",x"D0", -- 0x0190
    x"39",x"A5",x"59",x"DD",x"33",x"A2",x"D0",x"32", -- 0x0198
    x"20",x"E0",x"A1",x"CA",x"10",x"C0",x"A9",x"28", -- 0x01A0
    x"85",x"05",x"A9",x"3F",x"85",x"04",x"A9",x"A8", -- 0x01A8
    x"85",x"0A",x"A9",x"7C",x"85",x"09",x"20",x"21", -- 0x01B0
    x"A7",x"20",x"AC",x"A2",x"20",x"EE",x"A1",x"20", -- 0x01B8
    x"A7",x"A2",x"20",x"63",x"A6",x"20",x"2D",x"A4", -- 0x01C0
    x"20",x"84",x"A8",x"29",x"20",x"D0",x"ED",x"4C", -- 0x01C8
    x"07",x"A7",x"20",x"E0",x"A1",x"20",x"3B",x"A4", -- 0x01D0
    x"20",x"84",x"A8",x"29",x"20",x"D0",x"90",x"4C", -- 0x01D8
    x"07",x"A7",x"A5",x"48",x"85",x"04",x"A5",x"59", -- 0x01E0
    x"85",x"05",x"BD",x"6D",x"A2",x"4C",x"23",x"A0", -- 0x01E8
    x"A2",x"FF",x"A0",x"14",x"88",x"D0",x"FD",x"CA", -- 0x01F0
    x"D0",x"F8",x"60",x"20",x"28",x"30",x"38",x"48", -- 0x01F8
    x"50",x"58",x"60",x"68",x"70",x"78",x"80",x"40", -- 0x0200
    x"48",x"50",x"58",x"68",x"70",x"78",x"80",x"40", -- 0x0208
    x"48",x"50",x"58",x"60",x"68",x"70",x"78",x"80", -- 0x0210
    x"40",x"48",x"50",x"58",x"60",x"68",x"70",x"78", -- 0x0218
    x"80",x"48",x"50",x"58",x"60",x"10",x"18",x"20", -- 0x0220
    x"28",x"30",x"38",x"40",x"48",x"58",x"60",x"68", -- 0x0228
    x"70",x"78",x"80",x"88",x"90",x"70",x"70",x"70", -- 0x0230
    x"70",x"70",x"70",x"70",x"70",x"70",x"70",x"70", -- 0x0238
    x"70",x"78",x"78",x"78",x"78",x"78",x"78",x"78", -- 0x0240
    x"78",x"81",x"81",x"81",x"81",x"81",x"81",x"81", -- 0x0248
    x"81",x"81",x"89",x"89",x"89",x"89",x"89",x"89", -- 0x0250
    x"89",x"89",x"89",x"28",x"28",x"28",x"28",x"32", -- 0x0258
    x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"32", -- 0x0260
    x"32",x"32",x"32",x"32",x"32",x"32",x"32",x"59", -- 0x0268
    x"0F",x"15",x"12",x"45",x"0E",x"05",x"0D",x"09", -- 0x0270
    x"05",x"13",x"3A",x"45",x"16",x"09",x"0C",x"45", -- 0x0278
    x"19",x"05",x"13",x"57",x"0F",x"0C",x"17",x"0F", -- 0x0280
    x"0B",x"05",x"12",x"1A",x"4B",x"09",x"0C",x"0C", -- 0x0288
    x"05",x"12",x"02",x"0F",x"18",x"31",x"39",x"38", -- 0x0290
    x"32",x"43",x"12",x"05",x"01",x"14",x"09",x"16", -- 0x0298
    x"05",x"53",x"0F",x"06",x"14",x"17",x"01",x"12", -- 0x02A0
    x"05",x"20",x"AC",x"A2",x"E6",x"0C",x"A9",x"27", -- 0x02A8
    x"85",x"04",x"A9",x"78",x"85",x"05",x"20",x"3F", -- 0x02B0
    x"A9",x"A9",x"30",x"85",x"04",x"20",x"3F",x"A9", -- 0x02B8
    x"A9",x"2C",x"85",x"04",x"A9",x"81",x"85",x"05", -- 0x02C0
    x"20",x"8B",x"A9",x"A9",x"8B",x"85",x"05",x"4C", -- 0x02C8
    x"A6",x"A9",x"A5",x"E6",x"F8",x"18",x"69",x"01", -- 0x02D0
    x"85",x"E6",x"D8",x"29",x"0F",x"D0",x"08",x"A5", -- 0x02D8
    x"EA",x"C9",x"09",x"B0",x"02",x"E6",x"EA",x"20", -- 0x02E0
    x"07",x"A7",x"A5",x"E6",x"29",x"01",x"0A",x"AA", -- 0x02E8
    x"BD",x"FB",x"A2",x"85",x"00",x"BD",x"FC",x"A2", -- 0x02F0
    x"85",x"01",x"6C",x"00",x"00",x"14",x"A3",x"B8", -- 0x02F8
    x"A3",x"A2",x"FF",x"A9",x"14",x"E5",x"E6",x"29", -- 0x0300
    x"1F",x"69",x"01",x"85",x"F1",x"A4",x"F1",x"88", -- 0x0308
    x"D0",x"FD",x"CA",x"D0",x"F8",x"60",x"A9",x"64", -- 0x0310
    x"85",x"04",x"A9",x"58",x"85",x"05",x"20",x"5A", -- 0x0318
    x"A9",x"A9",x"05",x"85",x"F3",x"20",x"44",x"A3", -- 0x0320
    x"A9",x"96",x"8D",x"0A",x"90",x"A9",x"98",x"8D", -- 0x0328
    x"0B",x"90",x"20",x"FF",x"A2",x"20",x"44",x"A3", -- 0x0330
    x"E6",x"F3",x"A5",x"F3",x"C9",x"58",x"F0",x"2B", -- 0x0338
    x"20",x"44",x"A3",x"4C",x"30",x"A3",x"A9",x"58", -- 0x0340
    x"85",x"05",x"A5",x"F3",x"85",x"04",x"A9",x"A8", -- 0x0348
    x"85",x"0A",x"A9",x"54",x"85",x"09",x"20",x"21", -- 0x0350
    x"A7",x"A5",x"F3",x"18",x"69",x"08",x"85",x"04", -- 0x0358
    x"A9",x"A8",x"85",x"0A",x"A9",x"5C",x"85",x"09", -- 0x0360
    x"4C",x"21",x"A7",x"20",x"44",x"A3",x"20",x"C0", -- 0x0368
    x"AF",x"A9",x"64",x"85",x"F3",x"20",x"FF",x"A2", -- 0x0370
    x"A5",x"F3",x"85",x"04",x"20",x"5A",x"A9",x"E6", -- 0x0378
    x"F3",x"E6",x"0C",x"A5",x"F3",x"09",x"80",x"8D", -- 0x0380
    x"0D",x"90",x"C9",x"A0",x"F0",x"0A",x"A5",x"F3", -- 0x0388
    x"85",x"04",x"20",x"5A",x"A9",x"4C",x"73",x"A3", -- 0x0390
    x"A5",x"F3",x"85",x"04",x"A9",x"A8",x"85",x"0A", -- 0x0398
    x"A9",x"34",x"85",x"09",x"20",x"21",x"A7",x"A2", -- 0x03A0
    x"58",x"8A",x"48",x"20",x"FF",x"A2",x"20",x"9A", -- 0x03A8
    x"A8",x"8D",x"0D",x"90",x"68",x"AA",x"CA",x"D0", -- 0x03B0
    x"F0",x"60",x"A9",x"58",x"85",x"05",x"A9",x"05", -- 0x03B8
    x"85",x"F3",x"20",x"E6",x"A3",x"20",x"FF",x"A2", -- 0x03C0
    x"20",x"E6",x"A3",x"E6",x"F3",x"E6",x"0C",x"A5", -- 0x03C8
    x"0C",x"29",x"07",x"4A",x"09",x"C0",x"8D",x"0A", -- 0x03D0
    x"90",x"8D",x"0C",x"90",x"20",x"E6",x"A3",x"A5", -- 0x03D8
    x"F3",x"C9",x"9F",x"F0",x"14",x"4C",x"C3",x"A3", -- 0x03E0
    x"A5",x"F3",x"85",x"04",x"20",x"0F",x"A4",x"A5", -- 0x03E8
    x"F3",x"18",x"69",x"08",x"85",x"04",x"4C",x"5A", -- 0x03F0
    x"A9",x"A5",x"F3",x"18",x"69",x"08",x"85",x"04", -- 0x03F8
    x"20",x"5A",x"A9",x"A9",x"A8",x"85",x"0A",x"A9", -- 0x0400
    x"74",x"85",x"09",x"20",x"21",x"A7",x"4C",x"A5", -- 0x0408
    x"A3",x"A5",x"0C",x"4A",x"4A",x"29",x"01",x"F0", -- 0x0410
    x"0B",x"A9",x"A8",x"85",x"0A",x"A9",x"6C",x"85", -- 0x0418
    x"09",x"4C",x"21",x"A7",x"A9",x"A8",x"85",x"0A", -- 0x0420
    x"A9",x"64",x"85",x"09",x"4C",x"21",x"A7",x"8A", -- 0x0428
    x"48",x"A2",x"0F",x"20",x"3B",x"A4",x"CA",x"D0", -- 0x0430
    x"FA",x"68",x"AA",x"60",x"60",x"E6",x"0F",x"A5", -- 0x0438
    x"0F",x"29",x"3F",x"D0",x"F7",x"8A",x"48",x"A9", -- 0x0440
    x"A4",x"85",x"01",x"A9",x"7D",x"85",x"00",x"20", -- 0x0448
    x"7D",x"A0",x"20",x"7D",x"A0",x"20",x"7D",x"A0", -- 0x0450
    x"A0",x"00",x"B1",x"00",x"C9",x"FF",x"F0",x"14", -- 0x0458
    x"8D",x"0A",x"90",x"C8",x"B1",x"00",x"8D",x"0B", -- 0x0460
    x"90",x"C8",x"B1",x"00",x"8D",x"0C",x"90",x"E6", -- 0x0468
    x"0D",x"68",x"AA",x"60",x"A9",x"00",x"85",x"0D", -- 0x0470
    x"A9",x"FF",x"85",x"0F",x"4C",x"6F",x"A4",x"00", -- 0x0478
    x"E4",x"E4",x"00",x"E7",x"E7",x"00",x"E1",x"E1", -- 0x0480
    x"00",x"DB",x"DB",x"00",x"DB",x"DB",x"00",x"DF", -- 0x0488
    x"DF",x"00",x"D7",x"D7",x"00",x"D7",x"D7",x"00", -- 0x0490
    x"C9",x"C9",x"00",x"CF",x"CF",x"00",x"C3",x"C3", -- 0x0498
    x"00",x"B7",x"B7",x"00",x"B7",x"B7",x"00",x"BF", -- 0x04A0
    x"BF",x"00",x"AF",x"AF",x"00",x"AF",x"AF",x"C9", -- 0x04A8
    x"C9",x"00",x"CF",x"CF",x"00",x"C3",x"C3",x"00", -- 0x04B0
    x"B7",x"B7",x"00",x"B7",x"B7",x"00",x"BF",x"BF", -- 0x04B8
    x"00",x"B7",x"B7",x"00",x"B3",x"B3",x"00",x"AF", -- 0x04C0
    x"AF",x"00",x"AF",x"AF",x"00",x"00",x"00",x"00", -- 0x04C8
    x"00",x"00",x"00",x"EF",x"E4",x"EB",x"00",x"00", -- 0x04D0
    x"00",x"D7",x"BF",x"C9",x"D7",x"BF",x"CB",x"C3", -- 0x04D8
    x"00",x"CF",x"C3",x"00",x"E1",x"CF",x"D7",x"E1", -- 0x04E0
    x"CF",x"D7",x"CF",x"AF",x"AF",x"E1",x"AF",x"AF", -- 0x04E8
    x"E1",x"D7",x"C3",x"CF",x"D7",x"C3",x"E1",x"A3", -- 0x04F0
    x"A3",x"E1",x"A3",x"A3",x"E1",x"DB",x"C3",x"E1", -- 0x04F8
    x"DB",x"C3",x"E1",x"9F",x"9F",x"E1",x"9F",x"E1", -- 0x0500
    x"E1",x"D7",x"E4",x"E4",x"D7",x"E5",x"E5",x"AF", -- 0x0508
    x"E7",x"E7",x"AF",x"E1",x"E1",x"CF",x"E4",x"E4", -- 0x0510
    x"CF",x"E7",x"E7",x"AF",x"E7",x"E7",x"AF",x"DF", -- 0x0518
    x"DF",x"D7",x"E4",x"E4",x"D7",x"E4",x"E4",x"C3", -- 0x0520
    x"E1",x"E1",x"C3",x"E1",x"E1",x"E1",x"E1",x"E1", -- 0x0528
    x"00",x"E1",x"E1",x"E1",x"E1",x"E1",x"E1",x"E1", -- 0x0530
    x"E1",x"D7",x"BF",x"C9",x"D7",x"BF",x"CB",x"C3", -- 0x0538
    x"00",x"CF",x"C3",x"00",x"E1",x"CF",x"D7",x"E1", -- 0x0540
    x"CF",x"D7",x"CF",x"AF",x"AF",x"E1",x"AF",x"AF", -- 0x0548
    x"E1",x"D7",x"C3",x"CF",x"D7",x"C3",x"E1",x"A3", -- 0x0550
    x"A3",x"E1",x"A3",x"A3",x"E1",x"DB",x"C3",x"E1", -- 0x0558
    x"DB",x"C3",x"E1",x"9F",x"9F",x"E1",x"9F",x"9F", -- 0x0560
    x"E1",x"D4",x"DB",x"DB",x"D4",x"D7",x"D7",x"C9", -- 0x0568
    x"D4",x"D4",x"C9",x"DB",x"DB",x"DB",x"E1",x"E1", -- 0x0570
    x"DB",x"E7",x"E7",x"E4",x"E7",x"E7",x"E4",x"E4", -- 0x0578
    x"E4",x"E8",x"E1",x"E1",x"E8",x"DB",x"DB",x"EB", -- 0x0580
    x"E4",x"E4",x"EB",x"E4",x"E4",x"D7",x"E4",x"E4", -- 0x0588
    x"D7",x"E4",x"E4",x"DB",x"E4",x"E4",x"DB",x"E4", -- 0x0590
    x"E4",x"BF",x"BF",x"E4",x"BF",x"BF",x"E5",x"C3", -- 0x0598
    x"00",x"CF",x"C3",x"00",x"E1",x"CF",x"D7",x"E1", -- 0x05A0
    x"CF",x"D7",x"CF",x"AF",x"AF",x"E1",x"AF",x"AF", -- 0x05A8
    x"E1",x"D7",x"C3",x"CF",x"D7",x"C3",x"E1",x"A3", -- 0x05B0
    x"A3",x"E1",x"A3",x"A3",x"E1",x"DB",x"C3",x"E1", -- 0x05B8
    x"DB",x"C3",x"E1",x"9F",x"9F",x"E1",x"9F",x"E1", -- 0x05C0
    x"E1",x"D7",x"E4",x"E4",x"D7",x"E5",x"E5",x"AF", -- 0x05C8
    x"E7",x"E7",x"AF",x"E1",x"E1",x"CF",x"E4",x"E4", -- 0x05D0
    x"CF",x"E7",x"E7",x"AF",x"E7",x"E7",x"AF",x"E9", -- 0x05D8
    x"DF",x"D7",x"E4",x"E4",x"D7",x"E4",x"E4",x"C3", -- 0x05E0
    x"E1",x"E1",x"C3",x"E1",x"E1",x"E1",x"E1",x"E1", -- 0x05E8
    x"00",x"E1",x"E1",x"E1",x"E1",x"E1",x"E1",x"E1", -- 0x05F0
    x"E1",x"00",x"E1",x"E1",x"00",x"E4",x"E4",x"D7", -- 0x05F8
    x"E7",x"E7",x"D7",x"E1",x"E1",x"E7",x"E4",x"E4", -- 0x0600
    x"E7",x"E7",x"E7",x"DD",x"E7",x"E7",x"DD",x"E1", -- 0x0608
    x"E1",x"E1",x"E4",x"E4",x"E1",x"E1",x"E1",x"DB", -- 0x0610
    x"E7",x"E7",x"DB",x"E1",x"E1",x"E1",x"E4",x"E4", -- 0x0618
    x"E1",x"E7",x"E7",x"D9",x"E7",x"E7",x"D9",x"E1", -- 0x0620
    x"E1",x"E1",x"E4",x"E4",x"E1",x"E1",x"E1",x"D7", -- 0x0628
    x"E7",x"E7",x"D7",x"E1",x"E1",x"E7",x"E4",x"E4", -- 0x0630
    x"E7",x"E7",x"E7",x"AF",x"E7",x"E7",x"AF",x"DF", -- 0x0638
    x"DF",x"D7",x"E4",x"E4",x"E1",x"E7",x"E1",x"00", -- 0x0640
    x"E7",x"E1",x"D7",x"E7",x"E1",x"00",x"E7",x"E1", -- 0x0648
    x"C3",x"E7",x"E1",x"C3",x"E7",x"E1",x"C3",x"E7", -- 0x0650
    x"E1",x"C3",x"E7",x"E1",x"00",x"00",x"00",x"00", -- 0x0658
    x"00",x"00",x"FF",x"FF",x"FF",x"20",x"84",x"A8", -- 0x0660
    x"29",x"80",x"F0",x"13",x"A5",x"02",x"29",x"10", -- 0x0668
    x"F0",x"11",x"A5",x"02",x"29",x"08",x"F0",x"13", -- 0x0670
    x"A5",x"02",x"29",x"04",x"F0",x"09",x"60",x"EE", -- 0x0678
    x"00",x"90",x"60",x"CE",x"00",x"90",x"60",x"CE", -- 0x0680
    x"01",x"90",x"60",x"EE",x"01",x"90",x"60",x"A9", -- 0x0688
    x"8C",x"8D",x"05",x"90",x"A9",x"08",x"8D",x"0F", -- 0x0690
    x"90",x"A9",x"96",x"8D",x"02",x"90",x"A9",x"17", -- 0x0698
    x"8D",x"03",x"90",x"A9",x"0C",x"8D",x"00",x"90", -- 0x06A0
    x"A9",x"26",x"8D",x"01",x"90",x"A9",x"7F",x"8D", -- 0x06A8
    x"0E",x"90",x"A9",x"02",x"85",x"01",x"A9",x"00", -- 0x06B0
    x"85",x"00",x"A2",x"0B",x"A0",x"00",x"91",x"00", -- 0x06B8
    x"18",x"69",x"0B",x"C8",x"C0",x"16",x"D0",x"F6", -- 0x06C0
    x"48",x"A5",x"00",x"18",x"69",x"16",x"85",x"00", -- 0x06C8
    x"68",x"38",x"E9",x"F1",x"CA",x"D0",x"E5",x"A2", -- 0x06D0
    x"15",x"A9",x"07",x"9D",x"00",x"96",x"9D",x"DC", -- 0x06D8
    x"96",x"A9",x"06",x"9D",x"16",x"96",x"9D",x"C6", -- 0x06E0
    x"96",x"A9",x"02",x"9D",x"2C",x"96",x"9D",x"B0", -- 0x06E8
    x"96",x"A9",x"05",x"9D",x"42",x"96",x"9D",x"9A", -- 0x06F0
    x"96",x"A9",x"04",x"9D",x"58",x"96",x"9D",x"84", -- 0x06F8
    x"96",x"A9",x"03",x"9D",x"6E",x"96",x"CA",x"10", -- 0x0700
    x"D0",x"A9",x"00",x"85",x"00",x"A9",x"10",x"85", -- 0x0708
    x"01",x"A9",x"00",x"A8",x"91",x"00",x"E6",x"00", -- 0x0710
    x"D0",x"FA",x"E6",x"01",x"A5",x"01",x"C9",x"20", -- 0x0718
    x"D0",x"EF",x"60",x"8A",x"48",x"A5",x"04",x"4A", -- 0x0720
    x"4A",x"4A",x"AA",x"BD",x"70",x"A7",x"85",x"01", -- 0x0728
    x"BD",x"86",x"A7",x"18",x"65",x"05",x"85",x"00", -- 0x0730
    x"A5",x"01",x"69",x"00",x"85",x"01",x"A5",x"04", -- 0x0738
    x"29",x"07",x"85",x"0B",x"A0",x"07",x"B1",x"09", -- 0x0740
    x"85",x"13",x"A9",x"00",x"85",x"14",x"A6",x"0B", -- 0x0748
    x"F0",x"07",x"46",x"13",x"66",x"14",x"CA",x"D0", -- 0x0750
    x"F9",x"B1",x"00",x"45",x"13",x"91",x"00",x"98", -- 0x0758
    x"AA",x"09",x"B0",x"A8",x"B1",x"00",x"45",x"14", -- 0x0760
    x"91",x"00",x"8A",x"A8",x"88",x"10",x"D7",x"68", -- 0x0768
    x"AA",x"60",x"10",x"10",x"11",x"12",x"12",x"13", -- 0x0770
    x"14",x"14",x"15",x"16",x"16",x"17",x"18",x"18", -- 0x0778
    x"19",x"1A",x"1B",x"1B",x"1C",x"1D",x"1D",x"1E", -- 0x0780
    x"00",x"B0",x"60",x"10",x"C0",x"70",x"20",x"D0", -- 0x0788
    x"80",x"30",x"E0",x"90",x"40",x"F0",x"A0",x"50", -- 0x0790
    x"00",x"B0",x"60",x"10",x"C0",x"70",x"18",x"24", -- 0x0798
    x"42",x"CF",x"CF",x"42",x"24",x"18",x"18",x"2C", -- 0x07A0
    x"4E",x"C3",x"C3",x"42",x"24",x"18",x"18",x"3C", -- 0x07A8
    x"5A",x"C3",x"C3",x"42",x"24",x"18",x"18",x"34", -- 0x07B0
    x"72",x"C3",x"C3",x"42",x"24",x"18",x"18",x"24", -- 0x07B8
    x"42",x"E3",x"E3",x"42",x"24",x"18",x"18",x"24", -- 0x07C0
    x"42",x"C3",x"C3",x"72",x"34",x"18",x"18",x"24", -- 0x07C8
    x"42",x"C3",x"C3",x"5A",x"3C",x"18",x"18",x"24", -- 0x07D0
    x"42",x"C3",x"C3",x"4E",x"2C",x"18",x"30",x"30", -- 0x07D8
    x"11",x"7E",x"98",x"1C",x"16",x"34",x"18",x"18", -- 0x07E0
    x"90",x"7E",x"19",x"38",x"68",x"2C",x"24",x"42", -- 0x07E8
    x"A5",x"18",x"18",x"A5",x"42",x"24",x"30",x"62", -- 0x07F0
    x"13",x"1D",x"B8",x"C8",x"46",x"0C",x"3C",x"10", -- 0x07F8
    x"91",x"9F",x"F9",x"89",x"08",x"3C",x"0C",x"46", -- 0x0800
    x"C8",x"B8",x"1D",x"13",x"62",x"30",x"00",x"00", -- 0x0808
    x"18",x"34",x"34",x"18",x"00",x"00",x"00",x"00", -- 0x0810
    x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00", -- 0x0818
    x"3C",x"24",x"24",x"3C",x"00",x"00",x"00",x"7E", -- 0x0820
    x"42",x"42",x"42",x"42",x"7E",x"00",x"FF",x"81", -- 0x0828
    x"81",x"81",x"81",x"81",x"81",x"FF",x"10",x"10", -- 0x0830
    x"7C",x"10",x"10",x"10",x"38",x"7C",x"00",x"10", -- 0x0838
    x"10",x"36",x"50",x"10",x"38",x"7C",x"00",x"00", -- 0x0840
    x"10",x"10",x"14",x"52",x"B8",x"7C",x"00",x"00", -- 0x0848
    x"00",x"00",x"10",x"14",x"3A",x"7C",x"FF",x"80", -- 0x0850
    x"80",x"BC",x"C2",x"99",x"24",x"18",x"FC",x"1E", -- 0x0858
    x"1F",x"79",x"85",x"33",x"48",x"30",x"3C",x"7E", -- 0x0860
    x"F0",x"E0",x"E0",x"F0",x"7E",x"3C",x"3C",x"7E", -- 0x0868
    x"FF",x"F0",x"F0",x"FF",x"7E",x"3C",x"7E",x"C9", -- 0x0870
    x"ED",x"C9",x"FF",x"FF",x"FF",x"DB",x"3C",x"42", -- 0x0878
    x"BD",x"A5",x"A1",x"BD",x"42",x"3C",x"A9",x"7F", -- 0x0880
    x"8D",x"22",x"91",x"AD",x"20",x"91",x"29",x"80", -- 0x0888
    x"85",x"02",x"AD",x"1F",x"91",x"29",x"3C",x"05", -- 0x0890
    x"02",x"85",x"02",x"60",x"65",x"04",x"65",x"05", -- 0x0898
    x"6D",x"04",x"90",x"75",x"00",x"85",x"03",x"60", -- 0x08A0
    x"20",x"9A",x"A8",x"29",x"7F",x"69",x"14",x"60", -- 0x08A8
    x"A5",x"E6",x"49",x"FF",x"A8",x"88",x"D0",x"FD", -- 0x08B0
    x"60",x"FF",x"01",x"01",x"FF",x"FF",x"B5",x"15", -- 0x08B8
    x"F0",x"EE",x"C6",x"0C",x"20",x"37",x"A9",x"E6", -- 0x08C0
    x"0C",x"B5",x"37",x"A8",x"B5",x"15",x"18",x"79", -- 0x08C8
    x"B8",x"A8",x"95",x"15",x"B5",x"26",x"18",x"79", -- 0x08D0
    x"B7",x"A8",x"95",x"26",x"C9",x"A6",x"B0",x"2D", -- 0x08D8
    x"C9",x"02",x"90",x"29",x"B5",x"15",x"C9",x"A6", -- 0x08E0
    x"B0",x"31",x"C9",x"02",x"90",x"2D",x"A5",x"E7", -- 0x08E8
    x"F0",x"18",x"F5",x"15",x"69",x"03",x"C9",x"08", -- 0x08F0
    x"B0",x"10",x"A5",x"E8",x"F5",x"26",x"69",x"03", -- 0x08F8
    x"C9",x"08",x"B0",x"06",x"20",x"75",x"AE",x"95", -- 0x0900
    x"15",x"60",x"4C",x"37",x"A9",x"A9",x"FE",x"8D", -- 0x0908
    x"0C",x"90",x"B5",x"37",x"49",x"01",x"95",x"37", -- 0x0910
    x"4C",x"E2",x"A8",x"A9",x"FE",x"8D",x"0C",x"90", -- 0x0918
    x"B5",x"37",x"49",x"03",x"95",x"37",x"4C",x"EC", -- 0x0920
    x"A8",x"A7",x"A7",x"A7",x"A7",x"A7",x"A7",x"A7", -- 0x0928
    x"A7",x"9C",x"A4",x"AC",x"B4",x"BC",x"C4",x"CC", -- 0x0930
    x"D4",x"B5",x"15",x"85",x"04",x"B5",x"26",x"85", -- 0x0938
    x"05",x"A5",x"0C",x"4A",x"29",x"07",x"A8",x"B9", -- 0x0940
    x"27",x"A9",x"85",x"0A",x"B9",x"2F",x"A9",x"85", -- 0x0948
    x"09",x"4C",x"21",x"A7",x"A5",x"E1",x"85",x"04", -- 0x0950
    x"A5",x"E2",x"85",x"05",x"A5",x"0C",x"4A",x"4A", -- 0x0958
    x"4A",x"29",x"01",x"A8",x"B9",x"6F",x"A9",x"85", -- 0x0960
    x"0A",x"B9",x"71",x"A9",x"85",x"09",x"4C",x"21", -- 0x0968
    x"A7",x"A7",x"A7",x"DC",x"E4",x"A7",x"A7",x"A7", -- 0x0970
    x"A8",x"EC",x"F4",x"FC",x"04",x"A8",x"A8",x"A8", -- 0x0978
    x"A8",x"14",x"1C",x"24",x"2C",x"B5",x"48",x"85", -- 0x0980
    x"04",x"B5",x"59",x"85",x"05",x"A5",x"0C",x"4A", -- 0x0988
    x"29",x"03",x"A8",x"B9",x"73",x"A9",x"85",x"0A", -- 0x0990
    x"B9",x"77",x"A9",x"85",x"09",x"4C",x"21",x"A7", -- 0x0998
    x"A5",x"E3",x"85",x"04",x"A5",x"E4",x"85",x"05", -- 0x09A0
    x"A5",x"0C",x"4A",x"29",x"03",x"A8",x"B9",x"7B", -- 0x09A8
    x"A9",x"85",x"0A",x"B9",x"7F",x"A9",x"85",x"09", -- 0x09B0
    x"4C",x"21",x"A7",x"A5",x"E7",x"85",x"04",x"A5", -- 0x09B8
    x"E8",x"85",x"05",x"A9",x"A8",x"85",x"0A",x"A9", -- 0x09C0
    x"0C",x"85",x"09",x"4C",x"21",x"A7",x"A2",x"10", -- 0x09C8
    x"20",x"BC",x"A8",x"CA",x"10",x"FA",x"60",x"FF", -- 0x09D0
    x"01",x"01",x"FF",x"FF",x"A5",x"E3",x"F0",x"F6", -- 0x09D8
    x"C6",x"0C",x"20",x"9E",x"A9",x"E6",x"0C",x"A5", -- 0x09E0
    x"12",x"AA",x"A5",x"0C",x"3D",x"3B",x"AA",x"D0", -- 0x09E8
    x"05",x"20",x"DA",x"AF",x"85",x"11",x"A5",x"11", -- 0x09F0
    x"AA",x"A5",x"E3",x"18",x"7D",x"D6",x"A9",x"20", -- 0x09F8
    x"D3",x"AB",x"85",x"E3",x"A5",x"E4",x"18",x"7D", -- 0x0A00
    x"D5",x"A9",x"20",x"D3",x"AB",x"85",x"E4",x"A5", -- 0x0A08
    x"E7",x"F0",x"32",x"38",x"E5",x"E3",x"69",x"03", -- 0x0A10
    x"C9",x"08",x"B0",x"29",x"A5",x"E8",x"38",x"E5", -- 0x0A18
    x"E4",x"69",x"03",x"C9",x"08",x"B0",x"1E",x"20", -- 0x0A20
    x"75",x"AE",x"85",x"E3",x"60",x"04",x"00",x"05", -- 0x0A28
    x"07",x"09",x"00",x"10",x"10",x"00",x"04",x"05", -- 0x0A30
    x"07",x"09",x"10",x"00",x"10",x"7F",x"3F",x"1F", -- 0x0A38
    x"1F",x"0F",x"0F",x"07",x"07",x"4C",x"9E",x"A9", -- 0x0A40
    x"20",x"8B",x"A0",x"A9",x"03",x"85",x"EA",x"A9", -- 0x0A48
    x"00",x"85",x"EB",x"85",x"EC",x"85",x"ED",x"85", -- 0x0A50
    x"E6",x"20",x"07",x"A7",x"A2",x"10",x"A9",x"00", -- 0x0A58
    x"95",x"15",x"95",x"48",x"CA",x"10",x"F9",x"20", -- 0x0A60
    x"12",x"AB",x"BE",x"2B",x"AA",x"20",x"A6",x"A8", -- 0x0A68
    x"95",x"15",x"20",x"A6",x"A8",x"95",x"26",x"20", -- 0x0A70
    x"9A",x"A8",x"29",x"03",x"95",x"37",x"CA",x"10", -- 0x0A78
    x"EC",x"20",x"12",x"AB",x"BE",x"33",x"AA",x"20", -- 0x0A80
    x"A6",x"A8",x"95",x"48",x"20",x"A6",x"A8",x"95", -- 0x0A88
    x"59",x"20",x"9A",x"A8",x"29",x"07",x"95",x"6A", -- 0x0A90
    x"CA",x"10",x"EC",x"20",x"9E",x"AE",x"A2",x"13", -- 0x0A98
    x"A9",x"00",x"95",x"A3",x"CA",x"10",x"F9",x"A9", -- 0x0AA0
    x"00",x"85",x"E7",x"85",x"E5",x"85",x"E3",x"85", -- 0x0AA8
    x"10",x"85",x"0F",x"A9",x"02",x"85",x"E1",x"A9", -- 0x0AB0
    x"54",x"85",x"E2",x"20",x"52",x"A9",x"20",x"47", -- 0x0AB8
    x"A1",x"20",x"66",x"AD",x"20",x"77",x"AD",x"A9", -- 0x0AC0
    x"62",x"85",x"04",x"A9",x"08",x"85",x"05",x"A5", -- 0x0AC8
    x"E6",x"C9",x"10",x"90",x"06",x"20",x"47",x"AD", -- 0x0AD0
    x"4C",x"DC",x"AA",x"20",x"52",x"AD",x"E6",x"0C", -- 0x0AD8
    x"20",x"2C",x"AC",x"A5",x"0F",x"F0",x"25",x"A6", -- 0x0AE0
    x"0F",x"BD",x"CF",x"AF",x"8D",x"0D",x"90",x"C6", -- 0x0AE8
    x"0F",x"AD",x"0C",x"90",x"F0",x"03",x"EE",x"0C", -- 0x0AF0
    x"90",x"AD",x"0A",x"90",x"F0",x"03",x"CE",x"0A", -- 0x0AF8
    x"90",x"AD",x"0B",x"90",x"F0",x"03",x"CE",x"0B", -- 0x0B00
    x"90",x"4C",x"17",x"AE",x"A9",x"00",x"8D",x"0D", -- 0x0B08
    x"90",x"4C",x"EF",x"AA",x"A5",x"E6",x"29",x"07", -- 0x0B10
    x"A8",x"60",x"20",x"A9",x"AC",x"20",x"2A",x"AF", -- 0x0B18
    x"A5",x"0C",x"D0",x"0F",x"E6",x"10",x"A5",x"10", -- 0x0B20
    x"C9",x"03",x"D0",x"07",x"20",x"E6",x"AE",x"A9", -- 0x0B28
    x"00",x"85",x"10",x"20",x"60",x"AB",x"20",x"DA", -- 0x0B30
    x"A9",x"20",x"CC",x"A9",x"E6",x"0C",x"E6",x"0E", -- 0x0B38
    x"20",x"6D",x"AC",x"20",x"A9",x"AC",x"A2",x"10", -- 0x0B40
    x"B5",x"15",x"D0",x"94",x"B5",x"48",x"D0",x"90", -- 0x0B48
    x"CA",x"10",x"F5",x"20",x"0E",x"A1",x"20",x"D0", -- 0x0B50
    x"A2",x"20",x"07",x"A7",x"20",x"47",x"A1",x"4C", -- 0x0B58
    x"57",x"AA",x"A5",x"0C",x"29",x"1F",x"D0",x"0C", -- 0x0B60
    x"A2",x"10",x"20",x"9A",x"A8",x"29",x"07",x"95", -- 0x0B68
    x"6A",x"CA",x"10",x"F6",x"A2",x"10",x"B5",x"48", -- 0x0B70
    x"F0",x"4D",x"C6",x"0C",x"20",x"83",x"A9",x"E6", -- 0x0B78
    x"0C",x"B5",x"6A",x"A8",x"B5",x"48",x"18",x"79", -- 0x0B80
    x"CB",x"AB",x"95",x"48",x"B5",x"59",x"18",x"79", -- 0x0B88
    x"C9",x"AB",x"95",x"59",x"A5",x"59",x"B5",x"59", -- 0x0B90
    x"20",x"D3",x"AB",x"95",x"59",x"B5",x"48",x"20", -- 0x0B98
    x"D3",x"AB",x"95",x"48",x"A5",x"E7",x"F0",x"1C", -- 0x0BA0
    x"38",x"F5",x"48",x"69",x"03",x"C9",x"08",x"B0", -- 0x0BA8
    x"13",x"A5",x"E8",x"38",x"F5",x"59",x"69",x"03", -- 0x0BB0
    x"C9",x"08",x"B0",x"08",x"20",x"75",x"AE",x"95", -- 0x0BB8
    x"48",x"4C",x"C5",x"AB",x"20",x"83",x"A9",x"CA", -- 0x0BC0
    x"10",x"AC",x"60",x"FF",x"FF",x"00",x"01",x"01", -- 0x0BC8
    x"01",x"00",x"FF",x"FF",x"FF",x"C9",x"A8",x"B0", -- 0x0BD0
    x"05",x"C9",x"02",x"90",x"04",x"60",x"A9",x"A8", -- 0x0BD8
    x"60",x"A9",x"02",x"60",x"20",x"84",x"A8",x"49", -- 0x0BE0
    x"FF",x"29",x"9C",x"F0",x"20",x"C9",x"04",x"F0", -- 0x0BE8
    x"1F",x"C9",x"84",x"F0",x"1E",x"C9",x"80",x"F0", -- 0x0BF0
    x"1D",x"C9",x"88",x"F0",x"1C",x"C9",x"08",x"F0", -- 0x0BF8
    x"1B",x"C9",x"18",x"F0",x"1A",x"C9",x"10",x"F0", -- 0x0C00
    x"19",x"C9",x"14",x"F0",x"18",x"A9",x"80",x"60", -- 0x0C08
    x"A9",x"00",x"60",x"4C",x"CF",x"AD",x"A9",x"02", -- 0x0C10
    x"60",x"4C",x"08",x"AE",x"A9",x"04",x"60",x"4C", -- 0x0C18
    x"F3",x"AD",x"A9",x"06",x"60",x"4C",x"E4",x"AD", -- 0x0C20
    x"20",x"E2",x"AB",x"85",x"E5",x"60",x"20",x"26", -- 0x0C28
    x"AC",x"C6",x"0C",x"20",x"52",x"A9",x"E6",x"0C", -- 0x0C30
    x"A5",x"E5",x"C9",x"80",x"F0",x"23",x"AA",x"A5", -- 0x0C38
    x"E1",x"18",x"7D",x"CB",x"AB",x"20",x"D3",x"AB", -- 0x0C40
    x"C9",x"04",x"B0",x"02",x"A9",x"04",x"85",x"E1", -- 0x0C48
    x"A5",x"E2",x"18",x"7D",x"C9",x"AB",x"20",x"D3", -- 0x0C50
    x"AB",x"C9",x"04",x"B0",x"02",x"A9",x"04",x"85", -- 0x0C58
    x"E2",x"4C",x"52",x"A9",x"A5",x"0E",x"29",x"F0", -- 0x0C60
    x"F0",x"04",x"A9",x"00",x"85",x"0D",x"60",x"20", -- 0x0C68
    x"84",x"A8",x"29",x"20",x"D0",x"EE",x"20",x"26", -- 0x0C70
    x"AC",x"A5",x"E5",x"C9",x"80",x"F0",x"EF",x"A5", -- 0x0C78
    x"0D",x"D0",x"EB",x"A9",x"01",x"85",x"0D",x"85", -- 0x0C80
    x"0E",x"A5",x"E7",x"F0",x"03",x"20",x"B9",x"A9", -- 0x0C88
    x"A5",x"E1",x"85",x"E7",x"85",x"04",x"A5",x"E2", -- 0x0C90
    x"85",x"E8",x"85",x"05",x"A5",x"E5",x"85",x"E9", -- 0x0C98
    x"A9",x"8A",x"8D",x"0A",x"90",x"8D",x"0B",x"90", -- 0x0CA0
    x"4C",x"C1",x"A9",x"A5",x"E7",x"F0",x"BF",x"20", -- 0x0CA8
    x"B9",x"A9",x"A5",x"E9",x"AA",x"A5",x"E7",x"18", -- 0x0CB0
    x"7D",x"CB",x"AB",x"85",x"E7",x"A5",x"E8",x"18", -- 0x0CB8
    x"7D",x"C9",x"AB",x"85",x"E8",x"C9",x"A9",x"B0", -- 0x0CC0
    x"11",x"C9",x"02",x"90",x"0D",x"A5",x"E7",x"C9", -- 0x0CC8
    x"02",x"90",x"07",x"C9",x"A9",x"B0",x"03",x"4C", -- 0x0CD0
    x"B9",x"A9",x"A9",x"00",x"85",x"E7",x"60",x"4C", -- 0x0CD8
    x"46",x"AA",x"A2",x"FF",x"A9",x"8A",x"8D",x"0F", -- 0x0CE0
    x"90",x"A9",x"00",x"8D",x"0B",x"90",x"20",x"52", -- 0x0CE8
    x"A9",x"8E",x"0A",x"90",x"8E",x"0D",x"90",x"A0", -- 0x0CF0
    x"FF",x"A1",x"00",x"A1",x"00",x"A1",x"00",x"A1", -- 0x0CF8
    x"00",x"88",x"D0",x"F5",x"CA",x"D0",x"E7",x"A9", -- 0x0D00
    x"08",x"8D",x"0F",x"90",x"A5",x"EA",x"F0",x"CF", -- 0x0D08
    x"C6",x"EA",x"20",x"D1",x"AE",x"4C",x"99",x"AA", -- 0x0D10
    x"A0",x"00",x"B1",x"07",x"F0",x"19",x"C9",x"10", -- 0x0D18
    x"B0",x"06",x"20",x"52",x"AD",x"4C",x"2B",x"AD", -- 0x0D20
    x"B1",x"07",x"20",x"47",x"AD",x"C8",x"C0",x"03", -- 0x0D28
    x"D0",x"F6",x"A9",x"00",x"4C",x"52",x"AD",x"C8", -- 0x0D30
    x"C0",x"03",x"D0",x"DE",x"4C",x"30",x"AD",x"48", -- 0x0D38
    x"A5",x"04",x"18",x"69",x"08",x"85",x"04",x"68", -- 0x0D40
    x"60",x"85",x"F1",x"4A",x"4A",x"4A",x"4A",x"20", -- 0x0D48
    x"52",x"AD",x"A5",x"F1",x"29",x"0F",x"20",x"5B", -- 0x0D50
    x"AD",x"20",x"3D",x"AD",x"60",x"84",x"F2",x"18", -- 0x0D58
    x"69",x"30",x"20",x"23",x"A0",x"A4",x"F2",x"60", -- 0x0D60
    x"A9",x"00",x"85",x"04",x"85",x"05",x"A9",x"00", -- 0x0D68
    x"85",x"08",x"A9",x"EB",x"85",x"07",x"4C",x"16", -- 0x0D70
    x"AD",x"A9",x"62",x"85",x"04",x"A9",x"00",x"85", -- 0x0D78
    x"05",x"A9",x"00",x"85",x"08",x"A9",x"EE",x"85", -- 0x0D80
    x"07",x"4C",x"16",x"AD",x"8A",x"48",x"20",x"66", -- 0x0D88
    x"AD",x"20",x"77",x"AD",x"A5",x"ED",x"18",x"F8", -- 0x0D90
    x"69",x"05",x"85",x"ED",x"A5",x"EC",x"69",x"00", -- 0x0D98
    x"85",x"EC",x"A5",x"EB",x"69",x"00",x"85",x"EB", -- 0x0DA0
    x"D8",x"A5",x"EB",x"C5",x"EE",x"90",x"19",x"D0", -- 0x0DA8
    x"0E",x"A5",x"EC",x"C5",x"EF",x"90",x"11",x"D0", -- 0x0DB0
    x"06",x"A5",x"ED",x"C5",x"F0",x"90",x"09",x"A2", -- 0x0DB8
    x"02",x"B5",x"EB",x"95",x"EE",x"CA",x"10",x"F9", -- 0x0DC0
    x"20",x"77",x"AD",x"20",x"66",x"AD",x"68",x"AA", -- 0x0DC8
    x"60",x"A5",x"E1",x"C9",x"A7",x"B0",x"09",x"A5", -- 0x0DD0
    x"E2",x"C9",x"05",x"90",x"06",x"A9",x"01",x"60", -- 0x0DD8
    x"A9",x"00",x"60",x"A9",x"02",x"60",x"A5",x"E1", -- 0x0DE0
    x"C9",x"05",x"90",x"F4",x"A5",x"E2",x"C9",x"05", -- 0x0DE8
    x"90",x"12",x"A9",x"07",x"60",x"A5",x"E2",x"C9", -- 0x0DF0
    x"A7",x"B0",x"09",x"A5",x"E1",x"C9",x"05",x"90", -- 0x0DF8
    x"06",x"A9",x"05",x"60",x"A9",x"06",x"60",x"A9", -- 0x0E00
    x"04",x"60",x"A5",x"E2",x"C9",x"A7",x"B0",x"D3", -- 0x0E08
    x"A5",x"E1",x"C9",x"A7",x"B0",x"F1",x"A9",x"03", -- 0x0E10
    x"60",x"A2",x"10",x"B5",x"15",x"F0",x"19",x"A5", -- 0x0E18
    x"E1",x"38",x"F5",x"15",x"69",x"03",x"C9",x"08", -- 0x0E20
    x"B0",x"0E",x"A5",x"E2",x"38",x"F5",x"26",x"69", -- 0x0E28
    x"03",x"C9",x"08",x"B0",x"03",x"4C",x"E0",x"AC", -- 0x0E30
    x"B5",x"48",x"F0",x"19",x"A5",x"E1",x"38",x"F5", -- 0x0E38
    x"48",x"69",x"03",x"C9",x"08",x"B0",x"0E",x"A5", -- 0x0E40
    x"E2",x"38",x"F5",x"59",x"69",x"03",x"C9",x"08", -- 0x0E48
    x"B0",x"03",x"4C",x"E0",x"AC",x"CA",x"10",x"C3", -- 0x0E50
    x"A5",x"E3",x"F0",x"18",x"A5",x"E1",x"38",x"E5", -- 0x0E58
    x"E3",x"69",x"03",x"C9",x"08",x"B0",x"0D",x"A5", -- 0x0E60
    x"E2",x"E5",x"E4",x"69",x"03",x"E9",x"08",x"B0", -- 0x0E68
    x"03",x"4C",x"E0",x"AC",x"4C",x"18",x"AB",x"20", -- 0x0E70
    x"B9",x"A9",x"A5",x"E7",x"85",x"04",x"A5",x"E8", -- 0x0E78
    x"85",x"05",x"A9",x"A8",x"85",x"0A",x"A9",x"34", -- 0x0E80
    x"85",x"09",x"20",x"21",x"A7",x"8A",x"48",x"20", -- 0x0E88
    x"13",x"AF",x"68",x"AA",x"A9",x"09",x"85",x"0F", -- 0x0E90
    x"20",x"8A",x"AD",x"A9",x"00",x"85",x"E7",x"60", -- 0x0E98
    x"20",x"07",x"A7",x"A2",x"10",x"B5",x"15",x"F0", -- 0x0EA0
    x"09",x"85",x"04",x"B5",x"26",x"85",x"05",x"20", -- 0x0EA8
    x"3F",x"A9",x"CA",x"10",x"F0",x"A2",x"10",x"B5", -- 0x0EB0
    x"48",x"F0",x"09",x"85",x"04",x"B5",x"59",x"85", -- 0x0EB8
    x"05",x"20",x"8B",x"A9",x"CA",x"10",x"F0",x"60", -- 0x0EC0
    x"C9",x"14",x"B0",x"06",x"C9",x"00",x"F0",x"02", -- 0x0EC8
    x"69",x"14",x"60",x"A2",x"10",x"B5",x"15",x"20", -- 0x0ED0
    x"C6",x"AE",x"95",x"15",x"B5",x"48",x"20",x"C6", -- 0x0ED8
    x"AE",x"95",x"48",x"CA",x"10",x"EF",x"60",x"60", -- 0x0EE0
    x"A5",x"E3",x"D0",x"FB",x"20",x"9A",x"A8",x"29", -- 0x0EE8
    x"07",x"85",x"12",x"A5",x"E1",x"C9",x"58",x"90", -- 0x0EF0
    x"0B",x"20",x"DA",x"AF",x"85",x"11",x"A9",x"08", -- 0x0EF8
    x"20",x"04",x"AF",x"60",x"A9",x"A5",x"85",x"E3", -- 0x0F00
    x"20",x"A6",x"A8",x"85",x"E4",x"C6",x"0C",x"20", -- 0x0F08
    x"9E",x"A9",x"E6",x"0C",x"60",x"A2",x"13",x"B5", -- 0x0F10
    x"A3",x"F0",x"04",x"CA",x"10",x"F9",x"60",x"A5", -- 0x0F18
    x"E7",x"95",x"7B",x"A5",x"E8",x"95",x"8F",x"A9", -- 0x0F20
    x"05",x"95",x"A3",x"60",x"A5",x"0C",x"29",x"3F", -- 0x0F28
    x"D0",x"F9",x"A2",x"13",x"20",x"39",x"AF",x"CA", -- 0x0F30
    x"10",x"FA",x"60",x"B5",x"A3",x"F0",x"FB",x"C9", -- 0x0F38
    x"05",x"F0",x"14",x"C9",x"04",x"F0",x"0D",x"C9", -- 0x0F40
    x"03",x"F0",x"0F",x"C9",x"02",x"F0",x"11",x"C9", -- 0x0F48
    x"01",x"F0",x"13",x"60",x"20",x"6A",x"AF",x"D6", -- 0x0F50
    x"A3",x"60",x"20",x"70",x"AF",x"4C",x"55",x"AF", -- 0x0F58
    x"20",x"76",x"AF",x"4C",x"55",x"AF",x"20",x"7C", -- 0x0F60
    x"AF",x"4C",x"55",x"AF",x"20",x"88",x"AF",x"4C", -- 0x0F68
    x"96",x"AF",x"20",x"96",x"AF",x"4C",x"A4",x"AF", -- 0x0F70
    x"20",x"A4",x"AF",x"4C",x"B2",x"AF",x"4C",x"B2", -- 0x0F78
    x"AF",x"B5",x"7B",x"85",x"04",x"B5",x"8F",x"85", -- 0x0F80
    x"05",x"60",x"20",x"7F",x"AF",x"A9",x"A8",x"85", -- 0x0F88
    x"0A",x"A9",x"34",x"85",x"09",x"4C",x"21",x"A7", -- 0x0F90
    x"20",x"7F",x"AF",x"A9",x"A8",x"85",x"0A",x"A9", -- 0x0F98
    x"3C",x"85",x"09",x"4C",x"21",x"A7",x"20",x"7F", -- 0x0FA0
    x"AF",x"A9",x"A8",x"85",x"0A",x"A9",x"44",x"85", -- 0x0FA8
    x"09",x"4C",x"21",x"A7",x"20",x"7F",x"AF",x"A9", -- 0x0FB0
    x"A8",x"85",x"0A",x"A9",x"4C",x"85",x"09",x"4C", -- 0x0FB8
    x"21",x"A7",x"A9",x"00",x"8D",x"0A",x"90",x"8D", -- 0x0FC0
    x"0B",x"90",x"8D",x"0C",x"90",x"8D",x"0D",x"90", -- 0x0FC8
    x"60",x"99",x"81",x"9E",x"AC",x"C6",x"9B",x"C8", -- 0x0FD0
    x"B2",x"C6",x"BE",x"C9",x"A5",x"E3",x"C5",x"E1", -- 0x0FD8
    x"90",x"0C",x"A5",x"E4",x"C5",x"E2",x"90",x"03", -- 0x0FE0
    x"A9",x"03",x"60",x"A9",x"02",x"60",x"A5",x"E4", -- 0x0FE8
    x"C5",x"E2",x"90",x"03",x"A9",x"00",x"60",x"A9", -- 0x0FF0
    x"01",x"60",x"42",x"59",x"20",x"54",x"45",x"47", -- 0x0FF8
    x"52",x"32",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1000
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1008
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1010
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1018
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1020
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1028
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1030
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1038
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1040
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1048
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1050
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1058
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1060
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1068
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1070
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1078
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1080
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1088
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1090
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1098
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1100
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1108
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1110
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1118
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1120
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1128
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1130
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1138
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1140
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1148
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1150
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1158
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1160
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1168
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1170
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1178
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1180
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1188
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1190
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1198
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1200
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1208
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1210
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1218
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1220
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1228
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1230
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1238
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1240
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1248
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1250
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1258
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1260
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1268
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1270
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1278
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1280
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1288
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1290
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1298
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1300
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1308
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1310
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1318
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1320
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1328
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1330
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1338
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1340
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1348
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1350
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1358
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1360
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1368
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1370
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1378
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1380
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1388
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1390
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1398
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1400
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1408
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1410
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1418
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1420
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1428
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1430
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1438
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1440
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1448
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1450
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1458
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1460
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1468
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1470
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1478
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1480
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1488
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1490
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1498
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1500
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1508
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1510
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1518
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1520
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1528
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1530
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1538
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1540
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1548
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1550
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1558
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1560
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1568
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1570
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1578
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1580
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1588
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1590
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1598
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1600
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1608
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1610
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1618
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1620
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1628
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1630
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1638
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1640
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1648
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1650
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1658
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1660
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1668
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1670
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1678
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1680
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1688
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1690
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1698
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1700
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1708
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1710
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1718
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1720
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1728
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1730
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1738
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1740
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1748
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1750
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1758
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1760
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1768
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1770
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1778
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1780
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1788
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1790
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1798
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1800
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1808
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1810
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1818
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1820
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1828
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1830
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1838
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1840
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1848
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1850
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1858
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1860
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1868
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1870
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1878
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1880
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1888
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1890
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1898
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1900
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1908
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1910
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1918
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1920
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1928
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1930
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1938
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1940
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1948
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1950
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1958
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1960
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1968
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1970
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1978
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1980
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1988
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1990
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1998
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x1FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
     DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
