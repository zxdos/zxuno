library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library UNISIM;
use UNISIM.vcomponents.all;

entity vdp_vram_fill is
	port (
		cpu_clk	: in  STD_LOGIC;
		cpu_WE	: in  STD_LOGIC;
		cpu_A		: in  STD_LOGIC_VECTOR (13 downto 0);
		cpu_D_in	: in  STD_LOGIC_VECTOR (7 downto 0);
		cpu_D_out: out STD_LOGIC_VECTOR (7 downto 0);
		vdp_clk	: in  STD_LOGIC;
		vdp_A		: in  STD_LOGIC_VECTOR (13 downto 0);
		vdp_D_out: out STD_LOGIC_VECTOR (7 downto 0)
		);
end vdp_vram_fill;

architecture Behavioral of vdp_vram_fill is
begin
	RAMB16_S1_inst0 : RAMB16_S1_S1
	generic map (
    INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => X"000000000F000000000000000000000000000000000000000000000000000000",
    INIT_05 => X"0000000F000000000000000000000000000000000000F0000000000000000000",
    INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => X"0000000000000000000000000F00000000000000000000000000000F0F00000F",
    INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		CLKA => cpu_clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(0 downto 0),
		DOA => cpu_D_out(0 downto 0),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => not vdp_clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(0 downto 0),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst1 : RAMB16_S1_S1
	generic map (
    INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => X"000000000FF0F00000FF00F0000F00F0000F0F00000000000000000000000000",
    INIT_05 => X"000000FF000000000000F000000000000000F00000F0F0F00000000000000000",
    INIT_06 => X"00000FFF00FF000000FFF00F000F000000FF0FF00F000FF00000000000FFFFF0",
    INIT_07 => X"00000FF00000F000000F0F0000F000F00000000000000000000FFFF000FF0FF0",
    INIT_08 => X"0FFFF0F00000000F0F00000F000FFF000F00000F00FF0FF00FFFFFF0000FFFF0",
    INIT_09 => X"00FFFFF00FFFFFFF0FFFFFFF0F0000000F00000F00FFFFFF000000000FFFFFFF",
    INIT_0A => X"0FFFFFFF0000FFFF00FFFFFF0000000F00FF00F00FF00FF00F00000000000FF0",
    INIT_0B => X"0000000000000F00000000000FF00000000000000F00000F000000FF0FF000FF",
    INIT_0C => X"0FFFFF0000000000000FF0000FFFFFFF0000000000FFF0000FFFF00000000000",
    INIT_0D => X"00FFF0000FFFF0000FFFF000000000000F000F0000000000000000000FFFF000",
    INIT_0E => X"00FFFF00000FFF000FFFFF000000000000F000000000F000FFFFFF00000FF000",
    INIT_0F => X"00000000000000F00000000000000000000000000F000F00000FFF000F000F00",
    INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		CLKA => cpu_clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(1 downto 1),
		DOA => cpu_D_out(1 downto 1),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => not vdp_clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(1 downto 1),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst2 : RAMB16_S1_S1
	generic map (
    INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => X"0000000000FFF0F00F0F0FF000FFF0F00FFFFFFF000000FF0000000000000000",
    INIT_05 => X"00000FF0000000000000F000000000000000F00000FFFFF0000FFF000F00000F",
    INIT_06 => X"0000FFFF0FFFF00F0FFFFF0F0FFFFFFF0FFFFFFF0F00FFFF000000000FFFFFFF",
    INIT_07 => X"0000FFFF0000F000000F0F0000F000F0000000000000000000FFFFFF0FFFFFFF",
    INIT_08 => X"0FFFF0FF0000000F0F00000F00FFFFF00F00000F0FFFFFFF0FFFFFFF0F0F00FF",
    INIT_09 => X"0FFFFFFF0FFFFFFF0FFFFFFF0F0000000FF000FF0FFFFFFF0F00000F0FFFFFFF",
    INIT_0A => X"0FFFFFFF00FFFFFF0FFFFFFF0000000F0FFFF0FF0FFFFFFF0FFFFFF00000FFFF",
    INIT_0B => X"0F00000000000FF00FFFFFFF00FF00000F00000F0F0000FF00000FF000FF0FF0",
    INIT_0C => X"FFFFFF0000000F0F0F0FFF000FFFFFFF0F000F000FFFFF000FFFFF0000000F00",
    INIT_0D => X"0FFFFF000FFFFF000FFFFF000F0000000FF0FF000FFFFF0F0F0000000FFFFF00",
    INIT_0E => X"0FFFFF0000FFFF000FFFFF000F000F000FFF0F000000FF00FFFFFF0000FFFF00",
    INIT_0F => X"0000000000000FF00000F000000000000F00000F0F00FF0000FFFF000FF0FF00",
    INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		CLKA => cpu_clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(2 downto 2),
		DOA => cpu_D_out(2 downto 2),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => not vdp_clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(2 downto 2),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst3 : RAMB16_S1_S1
	generic map (
    INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => X"000000FF0FFF0FFF0FF0FF000FF0F0FF0FFFFFFF000000FF0F0FFFFF00000000",
    INIT_05 => X"0000FF000FF000000000F0000FF0000000FFFFF0000FFF0000FFFFF00FF000FF",
    INIT_06 => X"0FFFF00F0F00F00F0F000F0F0FFFFFFF0F00F00F0F0FF00F0FFFFFFF0F00FF0F",
    INIT_07 => X"0F0FF00F000F0F00000F0F00000F0F000FF00FF00FF00FF00FF0F00F0F00F00F",
    INIT_08 => X"0F00F00F0000F00F0F00F00F0FF000FF0F00000F0F00F00F0000F00F0F0FFF0F",
    INIT_09 => X"0F00000F000FF00000000FF00F00000000FF0FF00F0000000FFFFFFF0000F000",
    INIT_0A => X"00FF00000FFF00000F0000000FFFFFFF0F0FF00F000FF00F0FFFFFFF0000F00F",
    INIT_0B => X"0F000000000000FF0FFFFFFF000FF0000F00000F0F000FFF0FFFFF00000FFF00",
    INIT_0C => X"F0F00F0000000F0F0F0F0F000F000F000F000F000F000F000F0F0F0000000FFF",
    INIT_0D => X"0F000F0000000F000000FF000FFFFFFF00FFF000FFFFFF0F0FFFFF0F00000F00",
    INIT_0E => X"0FF000000FF000000F0000000F000F000F0F0F0000000F0000F00F0000F00F00",
    INIT_0F => X"0000000000000F0000FFFFF00FFFFFFF0FFF0FFF0F0FFF000FF0000000FFF000",
    INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		CLKA => cpu_clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(3 downto 3),
		DOA => cpu_D_out(3 downto 3),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => not vdp_clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(3 downto 3),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst4 : RAMB16_S1_S1
	generic map (
    INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => X"00000FFF0F0FF00F000FF0000FF0F0FF000F0F00000000000F0FFFFF00000000",
    INIT_05 => X"000FF0000FF000000000F000FFF0000000FFFFF0000FFF000FF000FF00FFFFF0",
    INIT_06 => X"0FFF000F0F00F0FF0F000F0F000F00FF0F00F00F0FFF000F0FFFFFFF0F0FF00F",
    INIT_07 => X"0F0F000F000F0F00000F0F00000F0F00FFF00FF00FF00FF00F00F00F0F00F00F",
    INIT_08 => X"0F00000F0000F00F0F00F00F0F00000F0FF000FF0F00F00F0000F00F0F0FFF0F",
    INIT_09 => X"0F00000F0000FF000000FF000F000000000FFF000F0000000FFFFFFF0000F000",
    INIT_0A => X"000FF0000FFF00000F0000000FFFFFFF0F00FF0F0000F00F0FF0000F0000F00F",
    INIT_0B => X"0F000000000000FF0F00000F0000FF000FFFFFFF0F00FF0F0FFFFF00000FFF00",
    INIT_0C => X"F0F00F000FFFFFFF0F0F0F000F000F000F000F000F000F000F0F0F00000000FF",
    INIT_0D => X"0F000F0000000F00000FF00000FFFFFF000F0000F000000000FFFF0F00000F00",
    INIT_0E => X"00FF00000FF000000F0000000FFFFFFF0F0F0F0000000F0000F00F0000F00F00",
    INIT_0F => X"0000000000000FF00FFF0FFF0FFFFFFF00FFFFF00FFF0F00FFF00000000F0000",
    INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		CLKA => cpu_clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(4 downto 4),
		DOA => cpu_D_out(4 downto 4),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => not vdp_clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(4 downto 4),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst5 : RAMB16_S1_S1
	generic map (
    INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => X"00000F000F00FFFF00FF0FF000F0FFF00FFFFFFF000000FF0000000000000000",
    INIT_05 => X"00FF0000000000000000F000F00000000000F00000FFFFF00F00000F000FFF00",
    INIT_06 => X"0000000F0FFFFFF00FF00FFF000F0FF00FF000FF0FF000FF00000FF00FFFFFFF",
    INIT_07 => X"000000FF00F000F0000F0F000000F000F0000000000000000F00FFFF0FFFFFFF",
    INIT_08 => X"0FFFFFFF0FFFFFFF0FFFFFFF0FFFFFFF00FFFFF00FFFFFFF0FFFFFFF0FF000FF",
    INIT_09 => X"0FFFFFFF00000FF000000FF00FFFFFFF0000F0000FF000000F00000F0FFFFFFF",
    INIT_0A => X"00FF000000FFFFFF0FFFFFFF0000000F0FF0FFFF0FFFFFFF0F00000F0FFFFFFF",
    INIT_0B => X"0F00000000000FF00F00000F00000FF00FFFFFFF0F0FF00F00000FF000FF0FF0",
    INIT_0C => X"F0FFFF000FFFFFF00FFFFF000FFFFF000FFFFF000FFFFFFF0FFF0F0000000000",
    INIT_0D => X"0FFFFF000FFFFF000000FF00000000000FFFFFFFF0000000000000000FFFFFFF",
    INIT_0E => X"0FF0000000FFFF000FFFFF0000FFFFFF0F0FFF000FFFFF0000FFFF00FFFFFF00",
    INIT_0F => X"00000000000000F00F00000F000000000000F0000FF00F00F0FFFF0000FFF000",
    INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		CLKA => cpu_clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(5 downto 5),
		DOA => cpu_D_out(5 downto 5),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => not vdp_clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(5 downto 5),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst6 : RAMB16_S1_S1
	generic map (
    INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => X"000000000FFFFFF00FF0F0F000F00F000FFFFFFF000000FF0000000000000000",
    INIT_05 => X"0FF00000000000000000F000000000000000F00000F0F0F00000000000000000",
    INIT_06 => X"0000000F00FFFF0000F00FFF000FFF0000F000F00F0000F000000F0000FFFFF0",
    INIT_07 => X"000000F000F000F0000F0F000000F000000000000000000000000FF000FF0FF0",
    INIT_08 => X"00FFFFF00FFFFFFF0FFFFFFF0FFFFFFF000FFF000FFFFFFF0FFFFFF000FFFFF0",
    INIT_09 => X"00FFFFF00FFFFFFF0FFFFFFF0FFFFFFF0FFFFFFF00F00000000000000FFFFFFF",
    INIT_0A => X"0FFFFFFF0000FFFF00FFFFFF0000000F00F00FF00FFFFFFF0FFFFFFF0FFFFFFF",
    INIT_0B => X"0F00000000000F0000000000000000FF000000000FFF000F000000FF0FF000FF",
    INIT_0C => X"000FF00000000F0000FFF00000FFF00000FFF0000FFFFFFF00F0000000000000",
    INIT_0D => X"00FFF0000FFFFF000FFFFF00000000000FFFFFFFF0000000000000000FFFFFFF",
    INIT_0E => X"0FFFFF00000FFF0000FFFF0000000F000F00F0000FFFFF00000FF000FFFFFF00",
    INIT_0F => X"0000000000000FF00000000000000000000000000F000F00000FFF000FF0FF00",
    INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		CLKA => cpu_clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(6 downto 6),
		DOA => cpu_D_out(6 downto 6),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => not vdp_clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(6 downto 6),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

	RAMB16_S1_inst7 : RAMB16_S1_S1
	generic map (
    INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => X"0000000000FF00000F00FF0000000000000F0F00000000000000000000000000",
    INIT_05 => X"0F000000000000000000000000000000000000000000F0000000000000000000",
    INIT_06 => X"000000000000000000000000000FF00000000000000000000000000000000000",
    INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => X"000000000FFFFFFF0FFFFFFF000000000FFFFFFF000000000000000000000000",
    INIT_0A => X"0FFFFFFF000000000000000000000000000000000000000000FFFFF000000000",
    INIT_0B => X"0F00000000000000000000000000000F000000000FF0000F0000000F0F00000F",
    INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => X"00000000000000000FFFFF000000000000000000000000000000000000000000",
    INIT_0E => X"00FFFF0000000000000000000000000000000000000000000000000000000000",
    INIT_0F => X"0000000000000F0000000000000000000000000000000000000000000F000F00",
    INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		CLKA => cpu_clk,
		ADDRA => cpu_A,
		DIA => cpu_D_in(7 downto 7),
		DOA => cpu_D_out(7 downto 7),
		ENA => '1',
		SSRA => '0',
		WEA => cpu_WE,

		CLKB => not vdp_clk,
		ADDRB => vdp_A,
		DIB => "0",
		DOB => vdp_D_out(7 downto 7),
		ENB => '1',
		SSRB => '0',
		WEB => '0'
	);

end Behavioral;

