-------------------------------------------------------------------------------
--
-- FPGA Colecovision
--
-- $Id: generic_ram.vhd,v 1.2 2006/01/05 23:31:32 arnim Exp $
--
-- Generic RTL flavour.
--
-- Characteristics of the synchronous RAM:
--   - memory is updated with rising clock edge
--   - no read-through-write capability
--
-------------------------------------------------------------------------------
--
-- Copyright (c) 2006, Arnim Laeuger (arnim.laeuger@gmx.net)
--
-- All rights reserved
--
-- Redistribution and use in source and synthezised forms, with or without
-- modification, are permitted provided that the following conditions are met:
--
-- Redistributions of source code must retain the above copyright notice,
-- this list of conditions and the following disclaimer.
--
-- Redistributions in synthesized form must reproduce the above copyright
-- notice, this list of conditions and the following disclaimer in the
-- documentation and/or other materials provided with the distribution.
--
-- Neither the name of the author nor the names of other contributors may
-- be used to endorse or promote products derived from this software without
-- specific prior written permission.
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
-- PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE
-- LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
-- CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
-- SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
-- INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
-- CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.
--
-- Please report bugs to the author, but before you do so, please
-- make sure that this is not a derivative work and that
-- you have the latest version of this file.
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity ram_init is

  generic (
    addr_width_g : integer := 13;
    data_width_g : integer := 8
  );
  port (
    clk_i : in  std_logic;
    a_i   : in  std_logic_vector(addr_width_g-1 downto 0);
    we_i  : in  std_logic;
    d_i   : in  std_logic_vector(data_width_g-1 downto 0);
    d_o   : out std_logic_vector(data_width_g-1 downto 0)
  );

end ram_init;


library ieee;
use ieee.numeric_std.all;

architecture rtl of ram_init is

  type mem_t is array (natural range 0 to 2**addr_width_g-1) of
    std_logic_vector(d_i'range);
  signal mem_q : mem_t := (
	 
	  x"31",x"26",x"3A",x"CD",x"0C",x"20",x"CD",x"BE", -- 0x0000
    x"22",x"C3",x"3F",x"20",x"21",x"D7",x"37",x"11", -- 0x0008
    x"B9",x"37",x"CD",x"35",x"20",x"11",x"B6",x"37", -- 0x0010
    x"21",x"54",x"37",x"01",x"51",x"37",x"CD",x"2A", -- 0x0018
    x"20",x"11",x"D7",x"37",x"21",x"B6",x"37",x"01", -- 0x0020
    x"B6",x"37",x"AF",x"ED",x"42",x"C5",x"4D",x"44", -- 0x0028
    x"E1",x"C8",x"ED",x"B0",x"C9",x"AF",x"E5",x"ED", -- 0x0030
    x"52",x"E1",x"C8",x"12",x"13",x"18",x"F7",x"00", -- 0x0038
    x"18",x"FE",x"04",x"05",x"C8",x"CB",x"3A",x"CB", -- 0x0040
    x"1B",x"10",x"FA",x"C9",x"F5",x"C5",x"E5",x"21", -- 0x0048
    x"00",x"00",x"CB",x"38",x"CB",x"19",x"38",x"0A", -- 0x0050
    x"78",x"B1",x"28",x"0D",x"CB",x"23",x"CB",x"12", -- 0x0058
    x"18",x"F0",x"19",x"CB",x"23",x"CB",x"12",x"18", -- 0x0060
    x"E9",x"EB",x"E1",x"C1",x"F1",x"C9",x"C5",x"E5", -- 0x0068
    x"F5",x"7C",x"EE",x"80",x"67",x"78",x"EE",x"80", -- 0x0070
    x"47",x"F1",x"A7",x"ED",x"42",x"E1",x"C1",x"C9", -- 0x0078
    x"B7",x"C8",x"FE",x"08",x"38",x"09",x"41",x"4C", -- 0x0080
    x"65",x"2E",x"00",x"D6",x"08",x"18",x"F2",x"29", -- 0x0088
    x"CB",x"11",x"CB",x"10",x"3D",x"20",x"F8",x"C9", -- 0x0090
    x"B7",x"C8",x"FE",x"08",x"38",x"09",x"6C",x"61", -- 0x0098
    x"48",x"06",x"00",x"D6",x"08",x"18",x"F2",x"CB", -- 0x00A0
    x"38",x"CB",x"19",x"CB",x"1C",x"CB",x"1D",x"3D", -- 0x00A8
    x"20",x"F5",x"C9",x"E3",x"D5",x"DD",x"E5",x"DD", -- 0x00B0
    x"21",x"00",x"00",x"DD",x"39",x"DD",x"56",x"09", -- 0x00B8
    x"DD",x"74",x"09",x"DD",x"5E",x"08",x"DD",x"75", -- 0x00C0
    x"08",x"D5",x"C5",x"F5",x"21",x"00",x"00",x"11", -- 0x00C8
    x"00",x"00",x"06",x"20",x"DD",x"4E",x"FD",x"DD", -- 0x00D0
    x"CB",x"FF",x"3E",x"DD",x"CB",x"FE",x"1E",x"DD", -- 0x00D8
    x"CB",x"07",x"1E",x"DD",x"CB",x"06",x"1E",x"30", -- 0x00E0
    x"12",x"7D",x"DD",x"86",x"04",x"6F",x"7C",x"DD", -- 0x00E8
    x"8E",x"05",x"67",x"7B",x"DD",x"8E",x"FC",x"5F", -- 0x00F0
    x"7A",x"89",x"57",x"DD",x"CB",x"04",x"26",x"DD", -- 0x00F8
    x"CB",x"05",x"16",x"DD",x"CB",x"FC",x"16",x"CB", -- 0x0100
    x"11",x"10",x"CC",x"DD",x"71",x"FD",x"42",x"4B", -- 0x0108
    x"F1",x"D1",x"D1",x"DD",x"E1",x"D1",x"33",x"33", -- 0x0110
    x"33",x"33",x"C9",x"EB",x"E3",x"F5",x"DD",x"E5", -- 0x0118
    x"DD",x"21",x"00",x"00",x"DD",x"39",x"C5",x"D5", -- 0x0120
    x"DD",x"56",x"09",x"DD",x"74",x"09",x"DD",x"5E", -- 0x0128
    x"08",x"DD",x"75",x"08",x"CD",x"43",x"21",x"E1", -- 0x0130
    x"C1",x"CD",x"DF",x"21",x"DD",x"E1",x"F1",x"D1", -- 0x0138
    x"33",x"33",x"C9",x"F5",x"21",x"00",x"00",x"01", -- 0x0140
    x"00",x"00",x"DD",x"36",x"F8",x"21",x"18",x"02", -- 0x0148
    x"19",x"37",x"DD",x"CB",x"FC",x"16",x"DD",x"CB", -- 0x0150
    x"FD",x"16",x"DD",x"CB",x"FE",x"16",x"DD",x"CB", -- 0x0158
    x"FF",x"16",x"DD",x"35",x"F8",x"28",x"2E",x"CB", -- 0x0160
    x"11",x"CB",x"10",x"CB",x"15",x"CB",x"14",x"ED", -- 0x0168
    x"52",x"38",x"DD",x"20",x"10",x"78",x"DD",x"96", -- 0x0170
    x"07",x"38",x"D5",x"20",x"08",x"79",x"DD",x"96", -- 0x0178
    x"06",x"38",x"CD",x"18",x"04",x"79",x"DD",x"96", -- 0x0180
    x"06",x"4F",x"78",x"DD",x"9E",x"07",x"47",x"30", -- 0x0188
    x"C1",x"2B",x"A7",x"18",x"BD",x"F1",x"E5",x"60", -- 0x0190
    x"69",x"C1",x"C9",x"EB",x"E3",x"F5",x"E5",x"21", -- 0x0198
    x"06",x"00",x"39",x"7E",x"A3",x"77",x"23",x"7E", -- 0x01A0
    x"A2",x"77",x"D1",x"23",x"7E",x"73",x"A1",x"4F", -- 0x01A8
    x"23",x"7E",x"72",x"A0",x"47",x"F1",x"D1",x"E1", -- 0x01B0
    x"C9",x"EB",x"E3",x"F5",x"E5",x"21",x"06",x"00", -- 0x01B8
    x"39",x"7E",x"B3",x"77",x"23",x"7E",x"B2",x"77", -- 0x01C0
    x"D1",x"23",x"7E",x"73",x"B1",x"4F",x"23",x"7E", -- 0x01C8
    x"72",x"B0",x"47",x"F1",x"D1",x"E1",x"C9",x"2C", -- 0x01D0
    x"C0",x"24",x"C0",x"0C",x"C0",x"04",x"C9",x"F5", -- 0x01D8
    x"7D",x"2F",x"6F",x"7C",x"2F",x"67",x"79",x"2F", -- 0x01E0
    x"4F",x"78",x"2F",x"47",x"F1",x"C9",x"C5",x"D5", -- 0x01E8
    x"5E",x"23",x"56",x"23",x"4E",x"23",x"46",x"EB", -- 0x01F0
    x"CD",x"B3",x"20",x"C3",x"FE",x"21",x"EB",x"70", -- 0x01F8
    x"2B",x"71",x"2B",x"72",x"2B",x"73",x"C9",x"F5", -- 0x0200
    x"7E",x"83",x"77",x"5F",x"23",x"7E",x"8A",x"77", -- 0x0208
    x"57",x"23",x"7E",x"89",x"77",x"4F",x"23",x"7E", -- 0x0210
    x"88",x"77",x"47",x"2B",x"2B",x"2B",x"F1",x"C9", -- 0x0218
    x"F5",x"7E",x"93",x"77",x"5F",x"23",x"7E",x"9A", -- 0x0220
    x"77",x"57",x"23",x"7E",x"99",x"77",x"4F",x"23", -- 0x0228
    x"7E",x"98",x"77",x"47",x"2B",x"2B",x"2B",x"F1", -- 0x0230
    x"C9",x"5E",x"23",x"56",x"23",x"4E",x"23",x"46", -- 0x0238
    x"EB",x"CD",x"80",x"20",x"C3",x"47",x"22",x"EB", -- 0x0240
    x"70",x"2B",x"71",x"2B",x"72",x"2B",x"73",x"C9", -- 0x0248
    x"E1",x"C5",x"D5",x"DD",x"E5",x"DD",x"21",x"00", -- 0x0250
    x"00",x"DD",x"39",x"E9",x"E1",x"C5",x"D5",x"DD", -- 0x0258
    x"E5",x"DD",x"21",x"00",x"00",x"DD",x"39",x"5E", -- 0x0260
    x"23",x"56",x"23",x"EB",x"39",x"F9",x"EB",x"E9", -- 0x0268
    x"DD",x"F9",x"DD",x"E1",x"D1",x"C1",x"C9",x"DD", -- 0x0270
    x"F9",x"DD",x"E1",x"D1",x"33",x"33",x"C9",x"F5", -- 0x0278
    x"E5",x"D5",x"C5",x"AF",x"EB",x"BE",x"ED",x"A0", -- 0x0280
    x"20",x"FB",x"C1",x"D1",x"E1",x"F1",x"C9",x"E5", -- 0x0288
    x"D5",x"C5",x"F5",x"AF",x"47",x"4F",x"ED",x"B1", -- 0x0290
    x"2B",x"EB",x"BE",x"ED",x"A0",x"20",x"FB",x"F1", -- 0x0298
    x"C1",x"D1",x"E1",x"C9",x"7E",x"BB",x"C8",x"B7", -- 0x02A0
    x"23",x"20",x"F9",x"21",x"00",x"00",x"C9",x"D5", -- 0x02A8
    x"21",x"54",x"37",x"E5",x"0E",x"12",x"1E",x"0C", -- 0x02B0
    x"CD",x"AD",x"36",x"E1",x"18",x"FE",x"CD",x"5C", -- 0x02B8
    x"22",x"A0",x"FF",x"FD",x"E5",x"CD",x"49",x"37", -- 0x02C0
    x"CD",x"41",x"37",x"CD",x"75",x"28",x"1E",x"00", -- 0x02C8
    x"CD",x"4A",x"25",x"1E",x"F4",x"CD",x"2F",x"37", -- 0x02D0
    x"CD",x"5C",x"25",x"CD",x"1F",x"37",x"3E",x"0B", -- 0x02D8
    x"01",x"24",x"00",x"ED",x"79",x"21",x"3E",x"00", -- 0x02E0
    x"39",x"EB",x"CD",x"67",x"2E",x"B7",x"28",x"04", -- 0x02E8
    x"5F",x"CD",x"AF",x"22",x"11",x"65",x"37",x"CD", -- 0x02F0
    x"A7",x"31",x"B7",x"28",x"04",x"5F",x"CD",x"AF", -- 0x02F8
    x"22",x"DD",x"70",x"A2",x"CD",x"3A",x"25",x"21", -- 0x0300
    x"6E",x"37",x"E5",x"0E",x"01",x"1E",x"0A",x"CD", -- 0x0308
    x"AD",x"36",x"E1",x"21",x"78",x"37",x"E5",x"0E", -- 0x0310
    x"02",x"1E",x"0A",x"CD",x"AD",x"36",x"E1",x"21", -- 0x0318
    x"82",x"37",x"E5",x"0E",x"03",x"59",x"CD",x"AD", -- 0x0320
    x"36",x"E1",x"DD",x"36",x"A3",x"00",x"21",x"0A", -- 0x0328
    x"00",x"39",x"E5",x"01",x"1B",x"00",x"11",x"B9", -- 0x0330
    x"37",x"CD",x"4B",x"32",x"E1",x"B7",x"20",x"2C", -- 0x0338
    x"DD",x"7E",x"A8",x"DD",x"B6",x"A9",x"28",x"24", -- 0x0340
    x"DD",x"34",x"A3",x"11",x"3B",x"00",x"21",x"B9", -- 0x0348
    x"37",x"CD",x"A4",x"22",x"72",x"21",x"B9",x"37", -- 0x0350
    x"E5",x"DD",x"7E",x"A3",x"C6",x"04",x"4F",x"1E", -- 0x0358
    x"04",x"CD",x"AD",x"36",x"E1",x"DD",x"7E",x"A3", -- 0x0360
    x"FE",x"0A",x"20",x"C2",x"21",x"B6",x"37",x"E5", -- 0x0368
    x"0E",x"05",x"CD",x"2C",x"25",x"E1",x"DD",x"36", -- 0x0370
    x"A1",x"05",x"DD",x"36",x"A4",x"00",x"1E",x"00", -- 0x0378
    x"CD",x"00",x"37",x"E5",x"FD",x"E1",x"CB",x"55", -- 0x0380
    x"28",x"2D",x"DD",x"4E",x"A3",x"06",x"00",x"21", -- 0x0388
    x"04",x"00",x"09",x"4D",x"44",x"DD",x"6E",x"A1", -- 0x0390
    x"26",x"00",x"CD",x"6E",x"20",x"30",x"18",x"21", -- 0x0398
    x"9E",x"37",x"E5",x"CD",x"29",x"25",x"E1",x"DD", -- 0x03A0
    x"34",x"A1",x"21",x"B6",x"37",x"E5",x"CD",x"29", -- 0x03A8
    x"25",x"E1",x"DD",x"34",x"A4",x"18",x"55",x"FD", -- 0x03B0
    x"E5",x"E1",x"CB",x"45",x"28",x"1F",x"3E",x"05", -- 0x03B8
    x"DD",x"BE",x"A1",x"30",x"18",x"21",x"9E",x"37", -- 0x03C0
    x"E5",x"CD",x"29",x"25",x"E1",x"DD",x"35",x"A1", -- 0x03C8
    x"21",x"B6",x"37",x"E5",x"CD",x"29",x"25",x"E1", -- 0x03D0
    x"DD",x"35",x"A4",x"18",x"2F",x"CB",x"5D",x"28", -- 0x03D8
    x"0B",x"AF",x"DD",x"B6",x"A2",x"28",x"0C",x"DD", -- 0x03E0
    x"35",x"A2",x"18",x"07",x"CB",x"4D",x"28",x"1C", -- 0x03E8
    x"DD",x"34",x"A2",x"DD",x"4E",x"A2",x"06",x"00", -- 0x03F0
    x"11",x"0E",x"01",x"CD",x"4C",x"20",x"7A",x"07", -- 0x03F8
    x"9F",x"4F",x"41",x"CD",x"38",x"34",x"DD",x"36", -- 0x0400
    x"A5",x"00",x"18",x"2F",x"FD",x"E5",x"E1",x"7C", -- 0x0408
    x"E6",x"C0",x"28",x"06",x"DD",x"36",x"A5",x"01", -- 0x0410
    x"18",x"21",x"DD",x"77",x"AA",x"DD",x"77",x"AB", -- 0x0418
    x"01",x"F0",x"0A",x"DD",x"6E",x"AA",x"DD",x"66", -- 0x0420
    x"AB",x"A7",x"ED",x"42",x"30",x"0A",x"DD",x"34", -- 0x0428
    x"AA",x"20",x"ED",x"DD",x"34",x"AB",x"18",x"E8", -- 0x0430
    x"C3",x"7E",x"23",x"AF",x"DD",x"B6",x"A5",x"CA", -- 0x0438
    x"04",x"23",x"FD",x"E5",x"E1",x"3E",x"40",x"AC", -- 0x0440
    x"B5",x"CA",x"1A",x"25",x"DD",x"4E",x"A4",x"06", -- 0x0448
    x"00",x"11",x"1B",x"00",x"CD",x"4C",x"20",x"D5", -- 0x0450
    x"DD",x"4E",x"A2",x"11",x"0E",x"01",x"CD",x"4C", -- 0x0458
    x"20",x"EB",x"D1",x"19",x"0E",x"11",x"09",x"EB", -- 0x0460
    x"7A",x"07",x"9F",x"4F",x"41",x"CD",x"38",x"34", -- 0x0468
    x"21",x"0A",x"00",x"39",x"E5",x"01",x"0D",x"00", -- 0x0470
    x"11",x"B9",x"37",x"CD",x"4B",x"32",x"E1",x"11", -- 0x0478
    x"0D",x"00",x"21",x"B9",x"37",x"CD",x"A4",x"22", -- 0x0480
    x"7D",x"B4",x"28",x"01",x"72",x"1E",x"20",x"21", -- 0x0488
    x"B9",x"37",x"CD",x"A4",x"22",x"7D",x"B4",x"28", -- 0x0490
    x"01",x"72",x"11",x"B9",x"37",x"21",x"14",x"00", -- 0x0498
    x"39",x"CD",x"7F",x"22",x"11",x"A1",x"37",x"21", -- 0x04A0
    x"14",x"00",x"39",x"CD",x"8F",x"22",x"21",x"A6", -- 0x04A8
    x"37",x"E5",x"0E",x"12",x"1E",x"04",x"CD",x"AD", -- 0x04B0
    x"36",x"E1",x"21",x"14",x"00",x"39",x"E5",x"0E", -- 0x04B8
    x"12",x"1E",x"0C",x"CD",x"AD",x"36",x"E1",x"11", -- 0x04C0
    x"AE",x"37",x"21",x"24",x"00",x"39",x"CD",x"7F", -- 0x04C8
    x"22",x"21",x"14",x"00",x"39",x"EB",x"21",x"24", -- 0x04D0
    x"00",x"39",x"CD",x"8F",x"22",x"EB",x"CD",x"A7", -- 0x04D8
    x"31",x"B7",x"28",x"04",x"5F",x"CD",x"AF",x"22", -- 0x04E0
    x"DD",x"36",x"B0",x"00",x"DD",x"36",x"B1",x"80", -- 0x04E8
    x"21",x"0A",x"00",x"39",x"E5",x"01",x"00",x"80", -- 0x04F0
    x"DD",x"5E",x"B0",x"DD",x"56",x"B1",x"CD",x"4B", -- 0x04F8
    x"32",x"E1",x"DD",x"77",x"A0",x"B7",x"20",x"08", -- 0x0500
    x"DD",x"7E",x"A8",x"DD",x"B6",x"A9",x"20",x"E0", -- 0x0508
    x"AF",x"DD",x"B6",x"A0",x"28",x"04",x"5F",x"CD", -- 0x0510
    x"AF",x"22",x"3E",x"04",x"D3",x"24",x"31",x"B9", -- 0x0518
    x"73",x"C3",x"6E",x"00",x"FD",x"E1",x"C3",x"70", -- 0x0520
    x"22",x"DD",x"4E",x"A1",x"1E",x"02",x"C3",x"AD", -- 0x0528
    x"36",x"CD",x"C0",x"08",x"2A",x"F6",x"73",x"19", -- 0x0530
    x"EB",x"C9",x"DD",x"E5",x"2A",x"F6",x"73",x"11", -- 0x0538
    x"00",x"03",x"3E",x"20",x"CD",x"82",x"1F",x"DD", -- 0x0540
    x"E1",x"C9",x"CD",x"50",x"22",x"DD",x"7E",x"02", -- 0x0548
    x"21",x"00",x"00",x"11",x"00",x"40",x"CD",x"82", -- 0x0550
    x"1F",x"C3",x"70",x"22",x"DD",x"E5",x"CD",x"7F", -- 0x0558
    x"1F",x"DD",x"E1",x"C9",x"CD",x"5C",x"22",x"00", -- 0x0560
    x"00",x"11",x"00",x"00",x"DD",x"4E",x"02",x"DD", -- 0x0568
    x"46",x"03",x"6B",x"62",x"A7",x"ED",x"42",x"30", -- 0x0570
    x"03",x"13",x"18",x"F0",x"C3",x"70",x"22",x"CD", -- 0x0578
    x"50",x"22",x"01",x"51",x"00",x"ED",x"59",x"C3", -- 0x0580
    x"70",x"22",x"C5",x"D5",x"3E",x"FF",x"01",x"51", -- 0x0588
    x"00",x"ED",x"79",x"0B",x"ED",x"50",x"7A",x"D1", -- 0x0590
    x"C1",x"C9",x"C5",x"DD",x"E5",x"D5",x"DD",x"E1", -- 0x0598
    x"3E",x"FF",x"01",x"51",x"00",x"ED",x"79",x"DD", -- 0x05A0
    x"2B",x"DD",x"E5",x"E1",x"7D",x"B4",x"20",x"F0", -- 0x05A8
    x"DD",x"E1",x"C1",x"C9",x"C5",x"CD",x"BA",x"25", -- 0x05B0
    x"C1",x"C9",x"3E",x"01",x"01",x"50",x"00",x"ED", -- 0x05B8
    x"79",x"C3",x"8A",x"25",x"CD",x"5C",x"22",x"FE", -- 0x05C0
    x"FF",x"DD",x"CB",x"02",x"7E",x"28",x"19",x"DD", -- 0x05C8
    x"CB",x"02",x"BE",x"21",x"00",x"00",x"E5",x"E5", -- 0x05D0
    x"1E",x"77",x"CD",x"C4",x"25",x"E1",x"E1",x"DD", -- 0x05D8
    x"77",x"FF",x"47",x"3E",x"01",x"B8",x"38",x"5B", -- 0x05E0
    x"CD",x"BA",x"25",x"AF",x"CD",x"BF",x"25",x"DD", -- 0x05E8
    x"5E",x"02",x"CD",x"7F",x"25",x"DD",x"4E",x"0A", -- 0x05F0
    x"DD",x"5E",x"0B",x"CD",x"7F",x"25",x"59",x"CD", -- 0x05F8
    x"7F",x"25",x"DD",x"5E",x"09",x"CD",x"7F",x"25", -- 0x0600
    x"DD",x"5E",x"08",x"CD",x"7F",x"25",x"DD",x"36", -- 0x0608
    x"FE",x"01",x"DD",x"7E",x"02",x"FE",x"40",x"20", -- 0x0610
    x"04",x"DD",x"36",x"FE",x"95",x"FE",x"48",x"20", -- 0x0618
    x"04",x"DD",x"36",x"FE",x"87",x"DD",x"5E",x"FE", -- 0x0620
    x"CD",x"7F",x"25",x"DD",x"36",x"FE",x"0A",x"CD", -- 0x0628
    x"8A",x"25",x"DD",x"77",x"FF",x"B7",x"F2",x"43", -- 0x0630
    x"26",x"DD",x"35",x"FE",x"DD",x"46",x"FE",x"04", -- 0x0638
    x"05",x"20",x"EC",x"DD",x"7E",x"FF",x"C3",x"70", -- 0x0640
    x"22",x"CD",x"5C",x"22",x"F6",x"FF",x"3E",x"01", -- 0x0648
    x"01",x"50",x"00",x"ED",x"79",x"11",x"64",x"00", -- 0x0650
    x"CD",x"9A",x"25",x"DD",x"70",x"F7",x"68",x"60", -- 0x0658
    x"E5",x"E5",x"1E",x"40",x"CD",x"C4",x"25",x"E1", -- 0x0660
    x"E1",x"3D",x"C2",x"6E",x"27",x"68",x"60",x"E5", -- 0x0668
    x"21",x"AA",x"01",x"E5",x"1E",x"48",x"CD",x"C4", -- 0x0670
    x"25",x"E1",x"E1",x"3D",x"C2",x"13",x"27",x"DD", -- 0x0678
    x"70",x"F6",x"DD",x"7E",x"F6",x"FE",x"04",x"30", -- 0x0680
    x"11",x"4F",x"21",x"04",x"00",x"39",x"09",x"E5", -- 0x0688
    x"CD",x"8A",x"25",x"E1",x"77",x"DD",x"34",x"F6", -- 0x0690
    x"18",x"E8",x"DD",x"46",x"FC",x"05",x"C2",x"6E", -- 0x0698
    x"27",x"DD",x"7E",x"FD",x"FE",x"AA",x"C2",x"6E", -- 0x06A0
    x"27",x"DD",x"36",x"F8",x"E8",x"DD",x"36",x"F9", -- 0x06A8
    x"03",x"DD",x"7E",x"F8",x"DD",x"B6",x"F9",x"28", -- 0x06B0
    x"15",x"21",x"00",x"40",x"E5",x"65",x"E5",x"1E", -- 0x06B8
    x"E9",x"CD",x"C4",x"25",x"E1",x"E1",x"B7",x"28", -- 0x06C0
    x"05",x"CD",x"84",x"27",x"18",x"E3",x"DD",x"7E", -- 0x06C8
    x"F8",x"DD",x"B6",x"F9",x"28",x"3B",x"21",x"00", -- 0x06D0
    x"00",x"E5",x"E5",x"1E",x"7A",x"CD",x"C4",x"25", -- 0x06D8
    x"E1",x"E1",x"B7",x"20",x"2C",x"DD",x"77",x"F6", -- 0x06E0
    x"DD",x"7E",x"F6",x"FE",x"04",x"30",x"13",x"4F", -- 0x06E8
    x"06",x"00",x"21",x"04",x"00",x"39",x"09",x"E5", -- 0x06F0
    x"CD",x"8A",x"25",x"E1",x"77",x"DD",x"34",x"F6", -- 0x06F8
    x"18",x"E6",x"DD",x"CB",x"FA",x"76",x"28",x"04", -- 0x0700
    x"3E",x"0C",x"18",x"02",x"3E",x"04",x"DD",x"77", -- 0x0708
    x"F7",x"18",x"5B",x"68",x"60",x"E5",x"E5",x"1E", -- 0x0710
    x"E9",x"CD",x"C4",x"25",x"E1",x"E1",x"47",x"3E", -- 0x0718
    x"01",x"B8",x"38",x"06",x"DD",x"36",x"F7",x"02", -- 0x0720
    x"18",x"03",x"DD",x"77",x"F7",x"DD",x"36",x"F8", -- 0x0728
    x"E8",x"DD",x"36",x"F9",x"03",x"DD",x"7E",x"F8", -- 0x0730
    x"DD",x"B6",x"F9",x"28",x"14",x"21",x"00",x"00", -- 0x0738
    x"E5",x"E5",x"1E",x"E9",x"CD",x"C4",x"25",x"E1", -- 0x0740
    x"E1",x"B7",x"28",x"05",x"CD",x"84",x"27",x"18", -- 0x0748
    x"E4",x"DD",x"7E",x"F8",x"DD",x"B6",x"F9",x"28", -- 0x0750
    x"11",x"21",x"00",x"00",x"E5",x"26",x"02",x"E5", -- 0x0758
    x"1E",x"50",x"CD",x"C4",x"25",x"E1",x"E1",x"B7", -- 0x0760
    x"28",x"04",x"DD",x"36",x"F7",x"00",x"DD",x"46", -- 0x0768
    x"F7",x"78",x"32",x"D4",x"37",x"CD",x"B4",x"25", -- 0x0770
    x"04",x"05",x"28",x"03",x"AF",x"18",x"02",x"3E", -- 0x0778
    x"01",x"C3",x"70",x"22",x"11",x"E8",x"03",x"CD", -- 0x0780
    x"64",x"25",x"DD",x"6E",x"F8",x"DD",x"66",x"F9", -- 0x0788
    x"2B",x"DD",x"75",x"F8",x"DD",x"74",x"F9",x"C9", -- 0x0790
    x"CD",x"5C",x"22",x"FC",x"FF",x"FD",x"E5",x"DD", -- 0x0798
    x"5E",x"0E",x"DD",x"56",x"0F",x"3A",x"D4",x"37", -- 0x07A0
    x"CB",x"5F",x"20",x"0B",x"D5",x"21",x"10",x"00", -- 0x07A8
    x"39",x"3E",x"09",x"CD",x"39",x"22",x"D1",x"DD", -- 0x07B0
    x"36",x"FD",x"01",x"D5",x"DD",x"6E",x"0A",x"DD", -- 0x07B8
    x"66",x"0B",x"E5",x"DD",x"6E",x"08",x"DD",x"66", -- 0x07C0
    x"09",x"E5",x"1E",x"51",x"CD",x"C4",x"25",x"E1", -- 0x07C8
    x"E1",x"B7",x"D1",x"C2",x"57",x"28",x"FD",x"21", -- 0x07D0
    x"E8",x"03",x"D5",x"11",x"64",x"00",x"CD",x"64", -- 0x07D8
    x"25",x"D1",x"CD",x"8A",x"25",x"DD",x"77",x"FC", -- 0x07E0
    x"3C",x"20",x"09",x"FD",x"2B",x"FD",x"E5",x"E1", -- 0x07E8
    x"7D",x"B4",x"20",x"E6",x"DD",x"46",x"FC",x"04", -- 0x07F0
    x"04",x"20",x"5C",x"DD",x"4E",x"0C",x"DD",x"46", -- 0x07F8
    x"0D",x"21",x"02",x"02",x"A7",x"ED",x"42",x"A7", -- 0x0800
    x"ED",x"52",x"DD",x"75",x"FE",x"DD",x"74",x"FF", -- 0x0808
    x"79",x"B0",x"28",x"0B",x"D5",x"DD",x"5E",x"0C", -- 0x0810
    x"DD",x"56",x"0D",x"CD",x"9A",x"25",x"D1",x"DD", -- 0x0818
    x"7E",x"02",x"DD",x"B6",x"03",x"28",x"1B",x"DD", -- 0x0820
    x"6E",x"02",x"DD",x"66",x"03",x"23",x"DD",x"75", -- 0x0828
    x"02",x"DD",x"74",x"03",x"2B",x"E5",x"CD",x"8A", -- 0x0830
    x"25",x"E1",x"77",x"1B",x"7B",x"B2",x"20",x"E7", -- 0x0838
    x"18",x"08",x"CD",x"8A",x"25",x"1B",x"7B",x"B2", -- 0x0840
    x"20",x"F8",x"DD",x"5E",x"FE",x"DD",x"56",x"FF", -- 0x0848
    x"CD",x"9A",x"25",x"DD",x"36",x"FD",x"00",x"CD", -- 0x0850
    x"B4",x"25",x"DD",x"7E",x"FD",x"FD",x"E1",x"C3", -- 0x0858
    x"70",x"22",x"DD",x"E5",x"3A",x"C4",x"73",x"F6", -- 0x0860
    x"20",x"4F",x"06",x"01",x"CD",x"D9",x"1F",x"CD", -- 0x0868
    x"DC",x"1F",x"DD",x"E1",x"C9",x"DD",x"E5",x"3A", -- 0x0870
    x"C4",x"73",x"E6",x"DF",x"4F",x"06",x"01",x"CD", -- 0x0878
    x"D9",x"1F",x"DD",x"E1",x"C9",x"CD",x"5C",x"22", -- 0x0880
    x"00",x"00",x"FD",x"E5",x"DD",x"5E",x"08",x"DD", -- 0x0888
    x"56",x"09",x"DD",x"6E",x"02",x"DD",x"66",x"03", -- 0x0890
    x"E5",x"FD",x"E1",x"7B",x"62",x"1B",x"B4",x"28", -- 0x0898
    x"0A",x"DD",x"46",x"04",x"FD",x"70",x"00",x"FD", -- 0x08A0
    x"23",x"18",x"F0",x"FD",x"E1",x"C3",x"70",x"22", -- 0x08A8
    x"CD",x"5C",x"22",x"FE",x"FF",x"FD",x"E5",x"DD", -- 0x08B0
    x"6E",x"02",x"DD",x"66",x"03",x"E5",x"FD",x"E1", -- 0x08B8
    x"59",x"50",x"AF",x"DD",x"77",x"FE",x"DD",x"77", -- 0x08C0
    x"FF",x"DD",x"6E",x"08",x"DD",x"66",x"09",x"2B", -- 0x08C8
    x"DD",x"75",x"08",x"DD",x"74",x"09",x"23",x"7D", -- 0x08D0
    x"B4",x"28",x"18",x"6B",x"62",x"13",x"4E",x"06", -- 0x08D8
    x"00",x"60",x"FD",x"6E",x"00",x"ED",x"42",x"DD", -- 0x08E0
    x"75",x"FE",x"DD",x"74",x"FF",x"7D",x"B4",x"FD", -- 0x08E8
    x"23",x"28",x"D6",x"DD",x"6E",x"FE",x"DD",x"66", -- 0x08F0
    x"FF",x"FD",x"E1",x"C3",x"70",x"22",x"CD",x"5C", -- 0x08F8
    x"22",x"FC",x"FF",x"FD",x"E5",x"FD",x"2A",x"D5", -- 0x0900
    x"37",x"01",x"02",x"00",x"DD",x"6E",x"02",x"DD", -- 0x0908
    x"66",x"03",x"A7",x"ED",x"42",x"38",x"56",x"FD", -- 0x0910
    x"4E",x"06",x"FD",x"46",x"07",x"DD",x"6E",x"02", -- 0x0918
    x"DD",x"66",x"03",x"ED",x"42",x"30",x"46",x"FD", -- 0x0920
    x"7E",x"00",x"FE",x"02",x"20",x"3F",x"21",x"02", -- 0x0928
    x"00",x"E5",x"DD",x"6E",x"02",x"29",x"E5",x"FD", -- 0x0930
    x"6E",x"0A",x"FD",x"66",x"0B",x"E5",x"FD",x"6E", -- 0x0938
    x"08",x"FD",x"66",x"09",x"E5",x"DD",x"6E",x"03", -- 0x0940
    x"26",x"00",x"5C",x"54",x"C1",x"09",x"EB",x"C1", -- 0x0948
    x"ED",x"4A",x"E5",x"D5",x"21",x"0A",x"00",x"39", -- 0x0950
    x"EB",x"CD",x"98",x"27",x"E1",x"E1",x"E1",x"E1", -- 0x0958
    x"B7",x"20",x"0A",x"DD",x"66",x"FD",x"DD",x"5E", -- 0x0960
    x"FC",x"B3",x"6F",x"18",x"03",x"21",x"01",x"00", -- 0x0968
    x"FD",x"E1",x"C3",x"70",x"22",x"FD",x"E5",x"DD", -- 0x0970
    x"E5",x"D5",x"FD",x"E1",x"DD",x"2A",x"D5",x"37", -- 0x0978
    x"21",x"06",x"00",x"ED",x"4B",x"D5",x"37",x"09", -- 0x0980
    x"46",x"23",x"66",x"68",x"01",x"FE",x"FF",x"09", -- 0x0988
    x"4D",x"44",x"FD",x"2B",x"FD",x"2B",x"FD",x"E5", -- 0x0990
    x"E1",x"A7",x"ED",x"42",x"38",x"07",x"01",x"00", -- 0x0998
    x"00",x"69",x"60",x"18",x"26",x"DD",x"6E",x"02", -- 0x09A0
    x"01",x"00",x"00",x"61",x"C5",x"E5",x"FD",x"E5", -- 0x09A8
    x"E1",x"CD",x"B3",x"20",x"C5",x"E5",x"DD",x"6E", -- 0x09B0
    x"10",x"DD",x"66",x"11",x"C1",x"09",x"EB",x"DD", -- 0x09B8
    x"6E",x"12",x"DD",x"66",x"13",x"C1",x"ED",x"4A", -- 0x09C0
    x"4D",x"44",x"EB",x"DD",x"E1",x"FD",x"E1",x"C9", -- 0x09C8
    x"C5",x"FD",x"E5",x"DD",x"E5",x"F5",x"D5",x"FD", -- 0x09D0
    x"E1",x"DD",x"2A",x"D5",x"37",x"EB",x"AF",x"77", -- 0x09D8
    x"23",x"77",x"6F",x"67",x"39",x"FD",x"4E",x"04", -- 0x09E0
    x"71",x"FD",x"46",x"05",x"23",x"70",x"3E",x"01", -- 0x09E8
    x"A9",x"B0",x"28",x"0F",x"DD",x"4E",x"06",x"DD", -- 0x09F0
    x"46",x"07",x"2B",x"56",x"23",x"66",x"6A",x"ED", -- 0x09F8
    x"42",x"38",x"04",x"3E",x"01",x"18",x"54",x"AF", -- 0x0A00
    x"28",x"19",x"6F",x"67",x"39",x"7A",x"23",x"B6", -- 0x0A08
    x"20",x"11",x"DD",x"7E",x"00",x"FE",x"03",x"20", -- 0x0A10
    x"0A",x"2B",x"DD",x"4E",x"0C",x"71",x"DD",x"46", -- 0x0A18
    x"0D",x"23",x"70",x"21",x"00",x"00",x"39",x"46", -- 0x0A20
    x"FD",x"70",x"06",x"23",x"66",x"FD",x"74",x"07", -- 0x0A28
    x"21",x"00",x"00",x"39",x"78",x"23",x"B6",x"28", -- 0x0A30
    x"09",x"2B",x"58",x"23",x"56",x"CD",x"75",x"29", -- 0x0A38
    x"18",x"0C",x"DD",x"4E",x"0E",x"DD",x"46",x"0F", -- 0x0A40
    x"DD",x"6E",x"0C",x"DD",x"66",x"0D",x"FD",x"75", -- 0x0A48
    x"08",x"FD",x"74",x"09",x"FD",x"71",x"0A",x"FD", -- 0x0A50
    x"70",x"0B",x"AF",x"E1",x"DD",x"E1",x"FD",x"E1", -- 0x0A58
    x"C1",x"C9",x"C5",x"FD",x"E5",x"DD",x"E5",x"F5", -- 0x0A60
    x"F5",x"D5",x"DD",x"E1",x"FD",x"2A",x"D5",x"37", -- 0x0A68
    x"21",x"00",x"00",x"39",x"1A",x"4F",x"13",x"1A", -- 0x0A70
    x"47",x"03",x"71",x"23",x"70",x"79",x"B0",x"28", -- 0x0A78
    x"49",x"DD",x"7E",x"08",x"DD",x"B6",x"09",x"DD", -- 0x0A80
    x"B6",x"0A",x"DD",x"B6",x"0B",x"28",x"3B",x"79", -- 0x0A88
    x"E6",x"0F",x"C2",x"40",x"2B",x"DD",x"6E",x"08", -- 0x0A90
    x"DD",x"66",x"09",x"DD",x"4E",x"0A",x"DD",x"46", -- 0x0A98
    x"0B",x"CD",x"D7",x"21",x"DD",x"75",x"08",x"DD", -- 0x0AA0
    x"74",x"09",x"DD",x"71",x"0A",x"DD",x"70",x"0B", -- 0x0AA8
    x"DD",x"7E",x"06",x"DD",x"B6",x"07",x"20",x"14", -- 0x0AB0
    x"FD",x"4E",x"04",x"FD",x"46",x"05",x"6F",x"67", -- 0x0AB8
    x"39",x"56",x"23",x"66",x"6A",x"A7",x"ED",x"42", -- 0x0AC0
    x"38",x"76",x"18",x"4D",x"06",x"04",x"21",x"00", -- 0x0AC8
    x"00",x"39",x"5E",x"23",x"56",x"CD",x"42",x"20", -- 0x0AD0
    x"FD",x"4E",x"02",x"06",x"00",x"0B",x"7B",x"A1", -- 0x0AD8
    x"67",x"7A",x"A0",x"B4",x"20",x"5A",x"21",x"02", -- 0x0AE0
    x"00",x"39",x"E5",x"DD",x"5E",x"06",x"DD",x"56", -- 0x0AE8
    x"07",x"CD",x"FE",x"28",x"4D",x"44",x"E1",x"71", -- 0x0AF0
    x"23",x"70",x"21",x"01",x"00",x"A7",x"ED",x"42", -- 0x0AF8
    x"38",x"04",x"3E",x"01",x"18",x"4B",x"FD",x"4E", -- 0x0B00
    x"06",x"FD",x"46",x"07",x"21",x"02",x"00",x"39", -- 0x0B08
    x"56",x"23",x"66",x"6A",x"A7",x"ED",x"42",x"38", -- 0x0B10
    x"04",x"3E",x"03",x"18",x"34",x"21",x"02",x"00", -- 0x0B18
    x"39",x"42",x"DD",x"70",x"06",x"23",x"66",x"DD", -- 0x0B20
    x"74",x"07",x"21",x"02",x"00",x"39",x"58",x"23", -- 0x0B28
    x"56",x"CD",x"75",x"29",x"DD",x"75",x"08",x"DD", -- 0x0B30
    x"74",x"09",x"DD",x"71",x"0A",x"DD",x"70",x"0B", -- 0x0B38
    x"21",x"00",x"00",x"39",x"46",x"23",x"66",x"68", -- 0x0B40
    x"E5",x"DD",x"E5",x"E1",x"C1",x"71",x"23",x"70", -- 0x0B48
    x"AF",x"E1",x"E1",x"DD",x"E1",x"FD",x"E1",x"C1", -- 0x0B50
    x"C9",x"FD",x"E5",x"DD",x"E5",x"F5",x"D5",x"DD", -- 0x0B58
    x"E1",x"C5",x"FD",x"E1",x"CD",x"D0",x"29",x"21", -- 0x0B60
    x"00",x"00",x"39",x"77",x"AF",x"B6",x"20",x"6A", -- 0x0B68
    x"21",x"20",x"00",x"E5",x"DD",x"7E",x"00",x"E6", -- 0x0B70
    x"0F",x"6F",x"29",x"29",x"29",x"29",x"29",x"E5", -- 0x0B78
    x"DD",x"6E",x"0A",x"DD",x"66",x"0B",x"E5",x"DD", -- 0x0B80
    x"6E",x"08",x"DD",x"66",x"09",x"E5",x"FD",x"E5", -- 0x0B88
    x"D1",x"CD",x"98",x"27",x"E1",x"E1",x"E1",x"E1", -- 0x0B90
    x"B7",x"28",x"02",x"3E",x"01",x"21",x"00",x"00", -- 0x0B98
    x"39",x"77",x"AF",x"B6",x"20",x"34",x"FD",x"46", -- 0x0BA0
    x"00",x"B0",x"20",x"04",x"36",x"03",x"18",x"2A", -- 0x0BA8
    x"FD",x"CB",x"0B",x"5E",x"20",x"15",x"21",x"0B", -- 0x0BB0
    x"00",x"E5",x"DD",x"4E",x"02",x"DD",x"46",x"03", -- 0x0BB8
    x"FD",x"E5",x"D1",x"CD",x"B0",x"28",x"F1",x"7D", -- 0x0BC0
    x"B4",x"28",x"0F",x"DD",x"E5",x"D1",x"CD",x"62", -- 0x0BC8
    x"2A",x"21",x"00",x"00",x"39",x"77",x"AF",x"B6", -- 0x0BD0
    x"28",x"96",x"21",x"00",x"00",x"39",x"7E",x"E1", -- 0x0BD8
    x"DD",x"E1",x"FD",x"E1",x"C9",x"CD",x"5C",x"22", -- 0x0BE0
    x"FA",x"FF",x"FD",x"E5",x"DD",x"6E",x"02",x"DD", -- 0x0BE8
    x"66",x"03",x"23",x"23",x"7E",x"23",x"66",x"6F", -- 0x0BF0
    x"E5",x"FD",x"E1",x"01",x"0B",x"00",x"C5",x"0E", -- 0x0BF8
    x"20",x"EB",x"CD",x"85",x"28",x"E1",x"DD",x"6E", -- 0x0C00
    x"04",x"DD",x"66",x"05",x"46",x"23",x"66",x"68", -- 0x0C08
    x"EB",x"DD",x"36",x"FB",x"00",x"DD",x"36",x"FC", -- 0x0C10
    x"00",x"DD",x"36",x"FD",x"08",x"DD",x"4E",x"FC", -- 0x0C18
    x"DD",x"34",x"FC",x"06",x"00",x"6B",x"62",x"09", -- 0x0C20
    x"46",x"DD",x"70",x"FA",x"3E",x"20",x"B8",x"30", -- 0x0C28
    x"05",x"78",x"FE",x"2F",x"20",x"03",x"C3",x"C2", -- 0x0C30
    x"2C",x"FE",x"2E",x"28",x"08",x"DD",x"7E",x"FB", -- 0x0C38
    x"DD",x"BE",x"FD",x"38",x"16",x"DD",x"7E",x"FD", -- 0x0C40
    x"FE",x"08",x"20",x"76",x"78",x"FE",x"2E",x"20", -- 0x0C48
    x"71",x"DD",x"36",x"FB",x"08",x"DD",x"36",x"FD", -- 0x0C50
    x"0B",x"18",x"C2",x"AF",x"28",x"3B",x"DD",x"4E", -- 0x0C58
    x"FD",x"47",x"0B",x"DD",x"6E",x"FB",x"67",x"CD", -- 0x0C60
    x"6E",x"20",x"30",x"2D",x"DD",x"4E",x"FC",x"DD", -- 0x0C68
    x"34",x"FC",x"44",x"6B",x"62",x"09",x"46",x"DD", -- 0x0C70
    x"70",x"FE",x"DD",x"4E",x"FB",x"DD",x"34",x"FB", -- 0x0C78
    x"47",x"FD",x"E5",x"E1",x"09",x"DD",x"46",x"FA", -- 0x0C80
    x"70",x"DD",x"4E",x"FB",x"DD",x"34",x"FB",x"47", -- 0x0C88
    x"FD",x"E5",x"E1",x"09",x"DD",x"46",x"FE",x"18", -- 0x0C90
    x"25",x"DD",x"7E",x"FA",x"FE",x"61",x"38",x"0F", -- 0x0C98
    x"3E",x"7A",x"DD",x"BE",x"FA",x"38",x"08",x"21", -- 0x0CA0
    x"02",x"00",x"39",x"7E",x"D6",x"20",x"77",x"DD", -- 0x0CA8
    x"4E",x"FB",x"DD",x"34",x"FB",x"06",x"00",x"FD", -- 0x0CB0
    x"E5",x"E1",x"09",x"DD",x"46",x"FA",x"70",x"C3", -- 0x0CB8
    x"1D",x"2C",x"DD",x"4E",x"FC",x"06",x"00",x"EB", -- 0x0CC0
    x"09",x"E5",x"DD",x"6E",x"04",x"DD",x"66",x"05", -- 0x0CC8
    x"C1",x"71",x"23",x"70",x"3E",x"20",x"DD",x"BE", -- 0x0CD0
    x"FA",x"38",x"04",x"3E",x"01",x"18",x"01",x"AF", -- 0x0CD8
    x"FD",x"77",x"0B",x"AF",x"FD",x"E1",x"C3",x"70", -- 0x0CE0
    x"22",x"CD",x"5C",x"22",x"FE",x"FF",x"FD",x"E5", -- 0x0CE8
    x"DD",x"6E",x"02",x"DD",x"66",x"03",x"E5",x"FD", -- 0x0CF0
    x"E1",x"DD",x"6E",x"08",x"DD",x"66",x"09",x"7E", -- 0x0CF8
    x"FE",x"20",x"20",x"0A",x"DD",x"34",x"08",x"20", -- 0x0D00
    x"F0",x"DD",x"34",x"09",x"18",x"EB",x"7E",x"FE", -- 0x0D08
    x"2F",x"20",x"08",x"DD",x"34",x"08",x"20",x"03", -- 0x0D10
    x"DD",x"34",x"09",x"AF",x"FD",x"77",x"04",x"FD", -- 0x0D18
    x"77",x"05",x"DD",x"6E",x"08",x"DD",x"66",x"09", -- 0x0D20
    x"3E",x"20",x"BE",x"38",x"13",x"FD",x"E5",x"D1", -- 0x0D28
    x"CD",x"D0",x"29",x"DD",x"77",x"FE",x"DD",x"6E", -- 0x0D30
    x"04",x"DD",x"66",x"05",x"36",x"00",x"18",x"6D", -- 0x0D38
    x"21",x"0C",x"00",x"39",x"4D",x"44",x"FD",x"E5", -- 0x0D40
    x"D1",x"CD",x"E5",x"2B",x"DD",x"77",x"FE",x"B7", -- 0x0D48
    x"20",x"5B",x"DD",x"4E",x"04",x"DD",x"46",x"05", -- 0x0D50
    x"FD",x"E5",x"D1",x"CD",x"59",x"2B",x"DD",x"77", -- 0x0D58
    x"FE",x"B7",x"28",x"14",x"FE",x"03",x"20",x"45", -- 0x0D60
    x"FD",x"6E",x"02",x"FD",x"66",x"03",x"01",x"0B", -- 0x0D68
    x"00",x"09",x"7E",x"B7",x"20",x"37",x"18",x"1B", -- 0x0D70
    x"FD",x"6E",x"02",x"FD",x"66",x"03",x"01",x"0B", -- 0x0D78
    x"00",x"09",x"7E",x"B7",x"20",x"27",x"69",x"60", -- 0x0D80
    x"DD",x"4E",x"04",x"DD",x"46",x"05",x"09",x"CB", -- 0x0D88
    x"66",x"20",x"06",x"DD",x"36",x"FE",x"04",x"18", -- 0x0D90
    x"14",x"21",x"1A",x"00",x"09",x"23",x"56",x"21", -- 0x0D98
    x"1A",x"00",x"09",x"4E",x"B1",x"FD",x"77",x"04", -- 0x0DA0
    x"FD",x"72",x"05",x"18",x"93",x"DD",x"7E",x"FE", -- 0x0DA8
    x"FD",x"E1",x"C3",x"70",x"22",x"C5",x"DD",x"E5", -- 0x0DB0
    x"D5",x"DD",x"E1",x"21",x"02",x"00",x"E5",x"21", -- 0x0DB8
    x"FE",x"01",x"E5",x"21",x"0A",x"00",x"39",x"4E", -- 0x0DC0
    x"23",x"46",x"23",x"5E",x"23",x"56",x"D5",x"C5", -- 0x0DC8
    x"DD",x"E5",x"D1",x"CD",x"98",x"27",x"E1",x"E1", -- 0x0DD0
    x"E1",x"E1",x"B7",x"28",x"05",x"3E",x"03",x"C3", -- 0x0DD8
    x"63",x"2E",x"DD",x"46",x"01",x"DD",x"5E",x"00", -- 0x0DE0
    x"B3",x"6F",x"78",x"B7",x"67",x"01",x"55",x"AA", -- 0x0DE8
    x"ED",x"42",x"28",x"04",x"3E",x"02",x"18",x"6B", -- 0x0DF0
    x"23",x"23",x"E5",x"2E",x"36",x"E5",x"2E",x"0A", -- 0x0DF8
    x"39",x"4E",x"23",x"46",x"23",x"5E",x"23",x"56", -- 0x0E00
    x"D5",x"C5",x"DD",x"E5",x"D1",x"CD",x"98",x"27", -- 0x0E08
    x"E1",x"E1",x"E1",x"E1",x"B7",x"20",x"12",x"DD", -- 0x0E10
    x"46",x"01",x"DD",x"5E",x"00",x"B3",x"6F",x"78", -- 0x0E18
    x"B7",x"67",x"01",x"46",x"41",x"ED",x"42",x"28", -- 0x0E20
    x"35",x"AF",x"28",x"35",x"21",x"02",x"00",x"E5", -- 0x0E28
    x"2E",x"52",x"E5",x"2E",x"0A",x"39",x"4E",x"23", -- 0x0E30
    x"46",x"23",x"5E",x"23",x"56",x"D5",x"C5",x"DD", -- 0x0E38
    x"E5",x"D1",x"CD",x"98",x"27",x"E1",x"E1",x"E1", -- 0x0E40
    x"E1",x"B7",x"20",x"15",x"DD",x"46",x"01",x"DD", -- 0x0E48
    x"5E",x"00",x"B3",x"6F",x"78",x"B7",x"67",x"01", -- 0x0E50
    x"46",x"41",x"ED",x"42",x"20",x"03",x"AF",x"18", -- 0x0E58
    x"02",x"3E",x"01",x"DD",x"E1",x"C1",x"C9",x"CD", -- 0x0E60
    x"5C",x"22",x"CA",x"FF",x"FD",x"E5",x"DD",x"6E", -- 0x0E68
    x"02",x"DD",x"66",x"03",x"E5",x"FD",x"E1",x"21", -- 0x0E70
    x"00",x"00",x"22",x"D5",x"37",x"FD",x"E5",x"E1", -- 0x0E78
    x"7D",x"B4",x"CA",x"88",x"31",x"CD",x"49",x"26", -- 0x0E80
    x"CB",x"47",x"28",x"05",x"3E",x"02",x"C3",x"89", -- 0x0E88
    x"31",x"21",x"00",x"00",x"E5",x"E5",x"2E",x"18", -- 0x0E90
    x"39",x"EB",x"CD",x"B5",x"2D",x"E1",x"E1",x"DD", -- 0x0E98
    x"77",x"CA",x"AF",x"DD",x"77",x"D0",x"DD",x"77", -- 0x0EA0
    x"D1",x"DD",x"77",x"D2",x"DD",x"77",x"D3",x"DD", -- 0x0EA8
    x"46",x"CA",x"05",x"20",x"67",x"21",x"10",x"00", -- 0x0EB0
    x"E5",x"21",x"BE",x"01",x"E5",x"6F",x"65",x"E5", -- 0x0EB8
    x"E5",x"2E",x"1C",x"39",x"EB",x"CD",x"98",x"27", -- 0x0EC0
    x"E1",x"E1",x"E1",x"E1",x"B7",x"28",x"06",x"DD", -- 0x0EC8
    x"36",x"CA",x"03",x"18",x"47",x"DD",x"7E",x"E0", -- 0x0ED0
    x"B7",x"28",x"41",x"DD",x"6E",x"E4",x"48",x"61", -- 0x0ED8
    x"C5",x"E5",x"DD",x"46",x"E5",x"4C",x"69",x"60", -- 0x0EE0
    x"41",x"C5",x"E5",x"DD",x"6E",x"E6",x"61",x"44", -- 0x0EE8
    x"4D",x"6C",x"C5",x"E5",x"DD",x"46",x"E7",x"6C", -- 0x0EF0
    x"CD",x"9B",x"31",x"CD",x"B9",x"21",x"CD",x"B9", -- 0x0EF8
    x"21",x"DD",x"75",x"D0",x"DD",x"74",x"D1",x"DD", -- 0x0F00
    x"71",x"D2",x"DD",x"70",x"D3",x"C5",x"E5",x"21", -- 0x0F08
    x"18",x"00",x"39",x"EB",x"CD",x"B5",x"2D",x"E1", -- 0x0F10
    x"E1",x"DD",x"77",x"CA",x"DD",x"7E",x"CA",x"FE", -- 0x0F18
    x"03",x"28",x"2B",x"AF",x"DD",x"B6",x"CA",x"C2", -- 0x0F20
    x"D8",x"30",x"21",x"24",x"00",x"E5",x"2E",x"0D", -- 0x0F28
    x"E5",x"DD",x"6E",x"D2",x"DD",x"66",x"D3",x"E5", -- 0x0F30
    x"DD",x"6E",x"D0",x"DD",x"66",x"D1",x"E5",x"21", -- 0x0F38
    x"1C",x"00",x"39",x"EB",x"CD",x"98",x"27",x"E1", -- 0x0F40
    x"E1",x"E1",x"E1",x"B7",x"28",x"05",x"3E",x"01", -- 0x0F48
    x"C3",x"89",x"31",x"DD",x"66",x"E6",x"4F",x"51", -- 0x0F50
    x"DD",x"5E",x"E5",x"79",x"B3",x"6F",x"DD",x"75", -- 0x0F58
    x"CC",x"41",x"DD",x"74",x"CD",x"DD",x"71",x"CE", -- 0x0F60
    x"DD",x"70",x"CF",x"7D",x"B4",x"20",x"2F",x"DD", -- 0x0F68
    x"6E",x"F3",x"61",x"C5",x"E5",x"DD",x"66",x"F4", -- 0x0F70
    x"4A",x"69",x"41",x"C5",x"E5",x"DD",x"6E",x"F5", -- 0x0F78
    x"61",x"44",x"4D",x"6A",x"C5",x"E5",x"DD",x"46", -- 0x0F80
    x"F6",x"CD",x"99",x"31",x"CD",x"B9",x"21",x"CD", -- 0x0F88
    x"B9",x"21",x"DD",x"75",x"CC",x"DD",x"74",x"CD", -- 0x0F90
    x"DD",x"71",x"CE",x"DD",x"70",x"CF",x"21",x"04", -- 0x0F98
    x"00",x"39",x"DD",x"5E",x"DF",x"4A",x"42",x"51", -- 0x0FA0
    x"CD",x"EE",x"21",x"DD",x"66",x"DE",x"0E",x"00", -- 0x0FA8
    x"79",x"DD",x"5E",x"DD",x"B3",x"6F",x"41",x"C5", -- 0x0FB0
    x"E5",x"DD",x"6E",x"D0",x"DD",x"66",x"D1",x"C1", -- 0x0FB8
    x"09",x"EB",x"DD",x"6E",x"D2",x"DD",x"66",x"D3", -- 0x0FC0
    x"C1",x"ED",x"4A",x"4D",x"44",x"EB",x"FD",x"75", -- 0x0FC8
    x"08",x"FD",x"74",x"09",x"FD",x"71",x"0A",x"FD", -- 0x0FD0
    x"70",x"0B",x"DD",x"46",x"DC",x"FD",x"70",x"02", -- 0x0FD8
    x"DD",x"66",x"E1",x"0E",x"00",x"51",x"DD",x"5E", -- 0x0FE0
    x"E0",x"79",x"B3",x"FD",x"77",x"04",x"FD",x"74", -- 0x0FE8
    x"05",x"DD",x"66",x"E3",x"4A",x"79",x"DD",x"5E", -- 0x0FF0
    x"E2",x"B3",x"6F",x"DD",x"75",x"D8",x"41",x"DD", -- 0x0FF8
    x"74",x"D9",x"DD",x"71",x"DA",x"DD",x"70",x"DB", -- 0x1000
    x"7D",x"B4",x"20",x"2F",x"DD",x"6E",x"EF",x"61", -- 0x1008
    x"C5",x"E5",x"DD",x"66",x"F0",x"4A",x"69",x"41", -- 0x1010
    x"C5",x"E5",x"DD",x"6E",x"F1",x"61",x"44",x"4D", -- 0x1018
    x"6A",x"C5",x"E5",x"DD",x"46",x"F2",x"CD",x"99", -- 0x1020
    x"31",x"CD",x"B9",x"21",x"CD",x"B9",x"21",x"DD", -- 0x1028
    x"75",x"D8",x"DD",x"74",x"D9",x"DD",x"71",x"DA", -- 0x1030
    x"DD",x"70",x"DB",x"FD",x"6E",x"02",x"4A",x"61", -- 0x1038
    x"42",x"C5",x"E5",x"CD",x"8E",x"31",x"D5",x"DD", -- 0x1040
    x"46",x"DE",x"4C",x"79",x"DD",x"6E",x"DD",x"B5", -- 0x1048
    x"5F",x"78",x"B7",x"57",x"69",x"ED",x"52",x"D1", -- 0x1050
    x"A7",x"ED",x"52",x"41",x"C5",x"E5",x"DD",x"6E", -- 0x1058
    x"D8",x"DD",x"66",x"D9",x"C1",x"09",x"EB",x"DD", -- 0x1060
    x"6E",x"DA",x"DD",x"66",x"DB",x"C1",x"ED",x"4A", -- 0x1068
    x"EB",x"A7",x"DD",x"4E",x"CC",x"DD",x"46",x"CD", -- 0x1070
    x"ED",x"42",x"EB",x"DD",x"4E",x"CE",x"DD",x"46", -- 0x1078
    x"CF",x"ED",x"42",x"CD",x"A1",x"31",x"C5",x"E5", -- 0x1080
    x"21",x"02",x"00",x"C1",x"09",x"EB",x"21",x"00", -- 0x1088
    x"00",x"C1",x"ED",x"4A",x"4D",x"44",x"EB",x"DD", -- 0x1090
    x"75",x"D4",x"DD",x"74",x"D5",x"DD",x"71",x"D6", -- 0x1098
    x"DD",x"70",x"D7",x"FD",x"75",x"06",x"FD",x"74", -- 0x10A0
    x"07",x"DD",x"36",x"CA",x"02",x"A7",x"01",x"F7", -- 0x10A8
    x"0F",x"ED",x"42",x"DD",x"6E",x"D6",x"DD",x"66", -- 0x10B0
    x"D7",x"01",x"00",x"00",x"ED",x"42",x"38",x"18", -- 0x10B8
    x"DD",x"6E",x"D4",x"DD",x"66",x"D5",x"01",x"F7", -- 0x10C0
    x"FF",x"ED",x"42",x"DD",x"6E",x"D6",x"DD",x"66", -- 0x10C8
    x"D7",x"01",x"00",x"00",x"ED",x"42",x"38",x"05", -- 0x10D0
    x"3E",x"07",x"C3",x"89",x"31",x"DD",x"46",x"CA", -- 0x10D8
    x"FD",x"70",x"00",x"AF",x"28",x"2D",x"78",x"FE", -- 0x10E0
    x"03",x"20",x"28",x"DD",x"6E",x"FB",x"41",x"61", -- 0x10E8
    x"C5",x"E5",x"DD",x"46",x"FC",x"4C",x"69",x"60", -- 0x10F0
    x"41",x"C5",x"E5",x"DD",x"6E",x"FD",x"61",x"44", -- 0x10F8
    x"4D",x"6C",x"C5",x"E5",x"DD",x"46",x"FE",x"6C", -- 0x1100
    x"CD",x"9B",x"31",x"CD",x"B9",x"21",x"CD",x"B9", -- 0x1108
    x"21",x"18",x"23",x"FD",x"6E",x"0A",x"FD",x"66", -- 0x1110
    x"0B",x"E5",x"FD",x"6E",x"08",x"FD",x"66",x"09", -- 0x1118
    x"E5",x"DD",x"6E",x"CC",x"DD",x"66",x"CD",x"C1", -- 0x1120
    x"09",x"EB",x"DD",x"6E",x"CE",x"DD",x"66",x"CF", -- 0x1128
    x"C1",x"ED",x"4A",x"4D",x"44",x"EB",x"FD",x"75", -- 0x1130
    x"0C",x"FD",x"74",x"0D",x"FD",x"71",x"0E",x"FD", -- 0x1138
    x"70",x"0F",x"CD",x"8E",x"31",x"EB",x"01",x"00", -- 0x1140
    x"00",x"C5",x"E5",x"FD",x"6E",x"08",x"FD",x"66", -- 0x1148
    x"09",x"C1",x"09",x"EB",x"FD",x"6E",x"0A",x"FD", -- 0x1150
    x"66",x"0B",x"C1",x"ED",x"4A",x"E5",x"D5",x"DD", -- 0x1158
    x"6E",x"CC",x"DD",x"66",x"CD",x"C1",x"09",x"EB", -- 0x1160
    x"DD",x"6E",x"CE",x"DD",x"66",x"CF",x"C1",x"ED", -- 0x1168
    x"4A",x"4D",x"44",x"EB",x"FD",x"75",x"10",x"FD", -- 0x1170
    x"74",x"11",x"FD",x"71",x"12",x"FD",x"70",x"13", -- 0x1178
    x"FD",x"36",x"01",x"00",x"FD",x"22",x"D5",x"37", -- 0x1180
    x"AF",x"FD",x"E1",x"C3",x"70",x"22",x"FD",x"5E", -- 0x1188
    x"04",x"FD",x"56",x"05",x"06",x"04",x"C3",x"42", -- 0x1190
    x"20",x"6A",x"65",x"4D",x"C3",x"B9",x"21",x"ED", -- 0x1198
    x"4A",x"4D",x"44",x"EB",x"C3",x"1B",x"21",x"CD", -- 0x11A0
    x"5C",x"22",x"C6",x"FF",x"FD",x"E5",x"FD",x"2A", -- 0x11A8
    x"D5",x"37",x"2A",x"D5",x"37",x"7D",x"B4",x"20", -- 0x11B0
    x"05",x"3E",x"06",x"C3",x"46",x"32",x"FD",x"36", -- 0x11B8
    x"01",x"00",x"21",x"30",x"00",x"39",x"DD",x"75", -- 0x11C0
    x"EA",x"DD",x"74",x"EB",x"DD",x"6E",x"02",x"DD", -- 0x11C8
    x"66",x"03",x"E5",x"21",x"06",x"00",x"39",x"4D", -- 0x11D0
    x"44",x"21",x"26",x"00",x"39",x"EB",x"CD",x"E9", -- 0x11D8
    x"2C",x"E1",x"B7",x"20",x"61",x"DD",x"B6",x"C8", -- 0x11E0
    x"28",x"06",x"DD",x"CB",x"D3",x"66",x"28",x"04", -- 0x11E8
    x"3E",x"03",x"18",x"52",x"DD",x"66",x"E3",x"0E", -- 0x11F0
    x"00",x"51",x"DD",x"5E",x"E2",x"79",x"B3",x"FD", -- 0x11F8
    x"77",x"1C",x"FD",x"74",x"1D",x"DD",x"6E",x"E4", -- 0x1200
    x"41",x"61",x"C5",x"E5",x"DD",x"66",x"E5",x"4A", -- 0x1208
    x"69",x"41",x"C5",x"E5",x"DD",x"6E",x"E6",x"61", -- 0x1210
    x"44",x"4D",x"6A",x"C5",x"E5",x"DD",x"46",x"E7", -- 0x1218
    x"CD",x"99",x"31",x"CD",x"B9",x"21",x"CD",x"B9", -- 0x1220
    x"21",x"FD",x"75",x"18",x"FD",x"74",x"19",x"FD", -- 0x1228
    x"71",x"1A",x"FD",x"70",x"1B",x"AF",x"FD",x"77", -- 0x1230
    x"14",x"FD",x"77",x"15",x"FD",x"77",x"16",x"FD", -- 0x1238
    x"77",x"17",x"FD",x"36",x"01",x"01",x"FD",x"E1", -- 0x1240
    x"C3",x"70",x"22",x"CD",x"5C",x"22",x"F0",x"FF", -- 0x1248
    x"FD",x"E5",x"DD",x"6E",x"02",x"DD",x"66",x"03", -- 0x1250
    x"DD",x"75",x"F2",x"DD",x"74",x"F3",x"FD",x"2A", -- 0x1258
    x"D5",x"37",x"DD",x"6E",x"08",x"DD",x"66",x"09", -- 0x1260
    x"AF",x"77",x"23",x"77",x"FD",x"E5",x"E1",x"7D", -- 0x1268
    x"B4",x"20",x"05",x"3E",x"06",x"C3",x"22",x"34", -- 0x1270
    x"FD",x"CB",x"01",x"46",x"20",x"05",x"3E",x"05", -- 0x1278
    x"C3",x"22",x"34",x"FD",x"6E",x"18",x"FD",x"66", -- 0x1280
    x"19",x"FD",x"4E",x"14",x"FD",x"46",x"15",x"ED", -- 0x1288
    x"42",x"EB",x"FD",x"6E",x"1A",x"FD",x"66",x"1B", -- 0x1290
    x"FD",x"4E",x"16",x"FD",x"46",x"17",x"ED",x"42", -- 0x1298
    x"4D",x"44",x"EB",x"DD",x"75",x"F4",x"DD",x"74", -- 0x12A0
    x"F5",x"DD",x"71",x"F6",x"DD",x"70",x"F7",x"DD", -- 0x12A8
    x"5E",x"04",x"DD",x"56",x"05",x"01",x"00",x"00", -- 0x12B0
    x"C5",x"D5",x"A7",x"C1",x"ED",x"42",x"DD",x"6E", -- 0x12B8
    x"F6",x"DD",x"66",x"F7",x"C1",x"ED",x"42",x"30", -- 0x12C0
    x"0C",x"DD",x"6E",x"F4",x"DD",x"66",x"F5",x"DD", -- 0x12C8
    x"75",x"04",x"DD",x"74",x"05",x"DD",x"7E",x"04", -- 0x12D0
    x"DD",x"B6",x"05",x"CA",x"22",x"34",x"FD",x"6E", -- 0x12D8
    x"14",x"FD",x"7E",x"15",x"E6",x"01",x"67",x"7D", -- 0x12E0
    x"B4",x"C2",x"70",x"33",x"CD",x"27",x"34",x"FD", -- 0x12E8
    x"7E",x"02",x"C6",x"FF",x"A5",x"DD",x"77",x"FE", -- 0x12F0
    x"20",x"30",x"FD",x"7E",x"14",x"FD",x"B6",x"15", -- 0x12F8
    x"FD",x"B6",x"16",x"FD",x"B6",x"17",x"20",x"08", -- 0x1300
    x"FD",x"6E",x"1C",x"FD",x"66",x"1D",x"18",x"09", -- 0x1308
    x"FD",x"5E",x"1E",x"FD",x"56",x"1F",x"CD",x"FE", -- 0x1310
    x"28",x"4D",x"44",x"21",x"01",x"00",x"A7",x"ED", -- 0x1318
    x"42",x"D2",x"1C",x"34",x"FD",x"71",x"1E",x"FD", -- 0x1320
    x"70",x"1F",x"FD",x"5E",x"1E",x"FD",x"56",x"1F", -- 0x1328
    x"CD",x"75",x"29",x"DD",x"75",x"F8",x"DD",x"74", -- 0x1330
    x"F9",x"DD",x"71",x"FA",x"DD",x"70",x"FB",x"7D", -- 0x1338
    x"B4",x"B1",x"B0",x"CA",x"1C",x"34",x"DD",x"6E", -- 0x1340
    x"FE",x"01",x"00",x"00",x"61",x"C5",x"E5",x"DD", -- 0x1348
    x"6E",x"F8",x"DD",x"66",x"F9",x"C1",x"09",x"EB", -- 0x1350
    x"DD",x"6E",x"FA",x"DD",x"66",x"FB",x"C1",x"ED", -- 0x1358
    x"4A",x"4D",x"44",x"EB",x"FD",x"75",x"20",x"FD", -- 0x1360
    x"74",x"21",x"FD",x"71",x"22",x"FD",x"70",x"23", -- 0x1368
    x"FD",x"4E",x"14",x"FD",x"7E",x"15",x"E6",x"01", -- 0x1370
    x"47",x"21",x"00",x"02",x"ED",x"42",x"DD",x"75", -- 0x1378
    x"F0",x"DD",x"74",x"F1",x"4D",x"44",x"DD",x"6E", -- 0x1380
    x"04",x"DD",x"66",x"05",x"A7",x"ED",x"42",x"30", -- 0x1388
    x"0C",x"DD",x"6E",x"04",x"DD",x"66",x"05",x"DD", -- 0x1390
    x"75",x"F0",x"DD",x"74",x"F1",x"DD",x"6E",x"F0", -- 0x1398
    x"DD",x"66",x"F1",x"E5",x"FD",x"6E",x"14",x"FD", -- 0x13A0
    x"7E",x"15",x"E6",x"01",x"67",x"E5",x"FD",x"6E", -- 0x13A8
    x"22",x"FD",x"66",x"23",x"E5",x"FD",x"6E",x"20", -- 0x13B0
    x"FD",x"66",x"21",x"E5",x"DD",x"7E",x"02",x"DD", -- 0x13B8
    x"B6",x"03",x"20",x"04",x"5F",x"57",x"18",x"06", -- 0x13C0
    x"DD",x"5E",x"F2",x"DD",x"56",x"F3",x"CD",x"98", -- 0x13C8
    x"27",x"E1",x"E1",x"E1",x"E1",x"B7",x"20",x"44", -- 0x13D0
    x"21",x"14",x"00",x"FD",x"E5",x"C1",x"09",x"DD", -- 0x13D8
    x"5E",x"F0",x"DD",x"56",x"F1",x"4F",x"47",x"CD", -- 0x13E0
    x"07",x"22",x"21",x"04",x"00",x"39",x"7E",x"DD", -- 0x13E8
    x"86",x"F0",x"77",x"23",x"7E",x"DD",x"8E",x"F1", -- 0x13F0
    x"77",x"21",x"16",x"00",x"39",x"7E",x"DD",x"96", -- 0x13F8
    x"F0",x"77",x"23",x"7E",x"DD",x"9E",x"F1",x"77", -- 0x1400
    x"DD",x"6E",x"08",x"DD",x"66",x"09",x"7E",x"DD", -- 0x1408
    x"86",x"F0",x"77",x"23",x"7E",x"DD",x"8E",x"F1", -- 0x1410
    x"77",x"C3",x"D5",x"32",x"FD",x"36",x"01",x"00", -- 0x1418
    x"3E",x"01",x"FD",x"E1",x"C3",x"70",x"22",x"FD", -- 0x1420
    x"4E",x"16",x"FD",x"46",x"17",x"FD",x"6E",x"14", -- 0x1428
    x"FD",x"66",x"15",x"3E",x"09",x"C3",x"98",x"20", -- 0x1430
    x"CD",x"5C",x"22",x"F2",x"FF",x"FD",x"E5",x"FD", -- 0x1438
    x"2A",x"D5",x"37",x"2A",x"D5",x"37",x"7D",x"B4", -- 0x1440
    x"20",x"05",x"3E",x"06",x"C3",x"A8",x"36",x"FD", -- 0x1448
    x"CB",x"01",x"46",x"20",x"05",x"3E",x"05",x"C3", -- 0x1450
    x"A8",x"36",x"FD",x"6E",x"18",x"FD",x"66",x"19", -- 0x1458
    x"DD",x"4E",x"02",x"DD",x"46",x"03",x"ED",x"42", -- 0x1460
    x"FD",x"6E",x"1A",x"FD",x"66",x"1B",x"DD",x"4E", -- 0x1468
    x"04",x"DD",x"46",x"05",x"ED",x"42",x"30",x"18", -- 0x1470
    x"FD",x"4E",x"1A",x"FD",x"46",x"1B",x"FD",x"6E", -- 0x1478
    x"18",x"DD",x"75",x"02",x"FD",x"66",x"19",x"DD", -- 0x1480
    x"74",x"03",x"DD",x"71",x"04",x"DD",x"70",x"05", -- 0x1488
    x"FD",x"4E",x"16",x"FD",x"46",x"17",x"FD",x"6E", -- 0x1490
    x"14",x"DD",x"75",x"F8",x"FD",x"66",x"15",x"DD", -- 0x1498
    x"74",x"F9",x"DD",x"71",x"FA",x"DD",x"70",x"FB", -- 0x14A0
    x"AF",x"FD",x"77",x"14",x"FD",x"77",x"15",x"FD", -- 0x14A8
    x"77",x"16",x"FD",x"77",x"17",x"DD",x"7E",x"02", -- 0x14B0
    x"DD",x"B6",x"03",x"DD",x"B6",x"04",x"DD",x"B6", -- 0x14B8
    x"05",x"CA",x"9F",x"36",x"FD",x"6E",x"02",x"01", -- 0x14C0
    x"00",x"00",x"61",x"3E",x"09",x"CD",x"80",x"20", -- 0x14C8
    x"DD",x"75",x"F4",x"DD",x"74",x"F5",x"DD",x"71", -- 0x14D0
    x"F6",x"DD",x"70",x"F7",x"DD",x"7E",x"F8",x"DD", -- 0x14D8
    x"B6",x"F9",x"DD",x"B6",x"FA",x"DD",x"B6",x"FB", -- 0x14E0
    x"CA",x"A2",x"35",x"C5",x"E5",x"21",x"FF",x"FF", -- 0x14E8
    x"E5",x"E5",x"DD",x"6E",x"F8",x"DD",x"66",x"F9", -- 0x14F0
    x"C1",x"09",x"EB",x"DD",x"6E",x"FA",x"DD",x"66", -- 0x14F8
    x"FB",x"C1",x"CD",x"9F",x"31",x"C5",x"E5",x"DD", -- 0x1500
    x"6E",x"F6",x"DD",x"66",x"F7",x"E5",x"DD",x"6E", -- 0x1508
    x"F4",x"DD",x"66",x"F5",x"E5",x"21",x"FF",x"FF", -- 0x1510
    x"E5",x"E5",x"DD",x"6E",x"02",x"DD",x"66",x"03", -- 0x1518
    x"C1",x"09",x"EB",x"DD",x"6E",x"04",x"DD",x"66", -- 0x1520
    x"05",x"C1",x"CD",x"9F",x"31",x"59",x"50",x"A7", -- 0x1528
    x"C1",x"ED",x"42",x"EB",x"C1",x"ED",x"42",x"38", -- 0x1530
    x"69",x"21",x"FF",x"FF",x"E5",x"E5",x"DD",x"6E", -- 0x1538
    x"F4",x"DD",x"66",x"F5",x"C1",x"09",x"EB",x"DD", -- 0x1540
    x"6E",x"F6",x"DD",x"66",x"F7",x"C1",x"ED",x"4A", -- 0x1548
    x"4D",x"44",x"EB",x"CD",x"DF",x"21",x"C5",x"E5", -- 0x1550
    x"21",x"FF",x"FF",x"E5",x"E5",x"DD",x"6E",x"F8", -- 0x1558
    x"DD",x"66",x"F9",x"C1",x"09",x"EB",x"DD",x"6E", -- 0x1560
    x"FA",x"DD",x"66",x"FB",x"C1",x"ED",x"4A",x"4D", -- 0x1568
    x"44",x"EB",x"CD",x"9B",x"21",x"FD",x"75",x"14", -- 0x1570
    x"FD",x"74",x"15",x"FD",x"71",x"16",x"FD",x"70", -- 0x1578
    x"17",x"21",x"12",x"00",x"39",x"FD",x"4E",x"16", -- 0x1580
    x"FD",x"46",x"17",x"FD",x"5E",x"14",x"FD",x"56", -- 0x1588
    x"15",x"CD",x"20",x"22",x"FD",x"6E",x"1E",x"DD", -- 0x1590
    x"75",x"F2",x"FD",x"66",x"1F",x"DD",x"74",x"F3", -- 0x1598
    x"18",x"12",x"FD",x"6E",x"1C",x"DD",x"75",x"F2", -- 0x15A0
    x"FD",x"66",x"1D",x"DD",x"74",x"F3",x"FD",x"75", -- 0x15A8
    x"1E",x"FD",x"74",x"1F",x"A7",x"DD",x"6E",x"F4", -- 0x15B0
    x"DD",x"66",x"F5",x"DD",x"4E",x"02",x"DD",x"46", -- 0x15B8
    x"03",x"ED",x"42",x"DD",x"6E",x"F6",x"DD",x"66", -- 0x15C0
    x"F7",x"DD",x"4E",x"04",x"DD",x"46",x"05",x"ED", -- 0x15C8
    x"42",x"30",x"65",x"DD",x"5E",x"F2",x"DD",x"56", -- 0x15D0
    x"F3",x"CD",x"FE",x"28",x"DD",x"75",x"F2",x"DD", -- 0x15D8
    x"74",x"F3",x"4D",x"44",x"21",x"01",x"00",x"A7", -- 0x15E0
    x"ED",x"42",x"30",x"11",x"FD",x"4E",x"06",x"FD", -- 0x15E8
    x"46",x"07",x"DD",x"6E",x"F2",x"DD",x"66",x"F3", -- 0x15F0
    x"A7",x"ED",x"42",x"38",x"03",x"C3",x"A2",x"36", -- 0x15F8
    x"DD",x"6E",x"F2",x"FD",x"75",x"1E",x"DD",x"66", -- 0x1600
    x"F3",x"FD",x"74",x"1F",x"21",x"14",x"00",x"FD", -- 0x1608
    x"E5",x"C1",x"09",x"DD",x"4E",x"F6",x"DD",x"46", -- 0x1610
    x"F7",x"DD",x"5E",x"F4",x"DD",x"56",x"F5",x"CD", -- 0x1618
    x"07",x"22",x"21",x"12",x"00",x"39",x"DD",x"4E", -- 0x1620
    x"F6",x"DD",x"46",x"F7",x"DD",x"5E",x"F4",x"DD", -- 0x1628
    x"56",x"F5",x"CD",x"20",x"22",x"C3",x"B4",x"35", -- 0x1630
    x"21",x"14",x"00",x"FD",x"E5",x"C1",x"09",x"DD", -- 0x1638
    x"4E",x"04",x"DD",x"46",x"05",x"DD",x"5E",x"02", -- 0x1640
    x"DD",x"56",x"03",x"CD",x"07",x"22",x"DD",x"5E", -- 0x1648
    x"F2",x"DD",x"56",x"F3",x"CD",x"75",x"29",x"DD", -- 0x1650
    x"75",x"FC",x"DD",x"74",x"FD",x"DD",x"71",x"FE", -- 0x1658
    x"DD",x"70",x"FF",x"7D",x"B4",x"B1",x"B0",x"28", -- 0x1660
    x"39",x"FD",x"6E",x"02",x"26",x"00",x"2B",x"7C", -- 0x1668
    x"07",x"9F",x"4F",x"41",x"C5",x"E5",x"CD",x"27", -- 0x1670
    x"34",x"CD",x"9B",x"21",x"C5",x"E5",x"DD",x"6E", -- 0x1678
    x"FC",x"DD",x"66",x"FD",x"C1",x"09",x"EB",x"DD", -- 0x1680
    x"6E",x"FE",x"DD",x"66",x"FF",x"C1",x"ED",x"4A", -- 0x1688
    x"4D",x"44",x"EB",x"FD",x"75",x"20",x"FD",x"74", -- 0x1690
    x"21",x"FD",x"71",x"22",x"FD",x"70",x"23",x"AF", -- 0x1698
    x"18",x"06",x"FD",x"36",x"01",x"00",x"3E",x"01", -- 0x16A0
    x"FD",x"E1",x"C3",x"70",x"22",x"CD",x"50",x"22", -- 0x16A8
    x"DD",x"56",x"04",x"DD",x"5E",x"02",x"CD",x"D4", -- 0x16B0
    x"36",x"D5",x"DD",x"5E",x"08",x"DD",x"56",x"09", -- 0x16B8
    x"CD",x"DD",x"36",x"06",x"00",x"4D",x"DD",x"6E", -- 0x16C0
    x"08",x"DD",x"66",x"09",x"D1",x"79",x"CD",x"DF", -- 0x16C8
    x"1F",x"C3",x"70",x"22",x"CD",x"C0",x"08",x"2A", -- 0x16D0
    x"F6",x"73",x"19",x"EB",x"C9",x"21",x"00",x"00", -- 0x16D8
    x"1A",x"B7",x"C8",x"23",x"13",x"18",x"F9",x"CD", -- 0x16E0
    x"50",x"22",x"51",x"CD",x"31",x"25",x"DD",x"6E", -- 0x16E8
    x"08",x"DD",x"66",x"09",x"DD",x"4E",x"0A",x"DD", -- 0x16F0
    x"46",x"0B",x"CD",x"DF",x"1F",x"C3",x"70",x"22", -- 0x16F8
    x"CD",x"50",x"22",x"CD",x"76",x"1F",x"DD",x"66", -- 0x1700
    x"02",x"2E",x"00",x"CD",x"79",x"1F",x"E5",x"DD", -- 0x1708
    x"66",x"02",x"2E",x"01",x"CD",x"79",x"1F",x"7C", -- 0x1710
    x"17",x"E1",x"B4",x"67",x"C3",x"70",x"22",x"DD", -- 0x1718
    x"E5",x"3A",x"C4",x"73",x"F6",x"40",x"4F",x"06", -- 0x1720
    x"01",x"CD",x"D9",x"1F",x"DD",x"E1",x"C9",x"CD", -- 0x1728
    x"50",x"22",x"DD",x"7E",x"02",x"21",x"00",x"20", -- 0x1730
    x"11",x"20",x"00",x"CD",x"82",x"1F",x"C3",x"70", -- 0x1738
    x"22",x"DD",x"E5",x"CD",x"85",x"1F",x"DD",x"E1", -- 0x1740
    x"C9",x"DD",x"E5",x"CD",x"E9",x"18",x"DD",x"E1", -- 0x1748
    x"C9",x"3D",x"3E",x"00",x"45",x"72",x"72",x"6F", -- 0x1750
    x"72",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x1758
    x"20",x"20",x"20",x"20",x"00",x"4D",x"45",x"4E", -- 0x1760
    x"55",x"2E",x"54",x"58",x"54",x"00",x"43",x"41", -- 0x1768
    x"52",x"54",x"20",x"4C",x"49",x"53",x"54",x"00", -- 0x1770
    x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D", -- 0x1778
    x"2D",x"00",x"52",x"2D",x"46",x"69",x"72",x"65", -- 0x1780
    x"3A",x"4C",x"6F",x"61",x"64",x"20",x"20",x"4C", -- 0x1788
    x"2D",x"46",x"69",x"72",x"65",x"3A",x"52",x"65", -- 0x1790
    x"73",x"74",x"61",x"72",x"74",x"00",x"20",x"20", -- 0x1798
    x"00",x"2E",x"72",x"6F",x"6D",x"00",x"4C",x"6F", -- 0x17A0
    x"61",x"64",x"69",x"6E",x"67",x"00",x"43",x"6F", -- 0x17A8
    x"6C",x"65",x"63",x"6F",x"2F",x"00",x"00",x"00", -- 0x17B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1800
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1808
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1810
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1818
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1820
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1828
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1830
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1838
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1840
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1848
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1850
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1858
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1860
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1868
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1870
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1878
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1880
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1888
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1890
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1898
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1900
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1908
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1910
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1918
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1920
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1928
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1930
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1938
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1940
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1948
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1950
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1958
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1960
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1968
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1970
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1978
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1980
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1988
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1990
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1998
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x1FF8
	 );


    -- pragma translate_off
    -- := (others => (others => '0'))
    -- pragma translate_on
   

begin

  mem: process (clk_i)
  begin

    if clk_i'event and clk_i = '1' then
      if we_i = '1' then
        mem_q(to_integer(unsigned(a_i))) <= d_i;
      end if;

      d_o <= mem_q(to_integer(unsigned(a_i)));
    end if;

  end process mem;

end rtl;
