-------------------------------------------------------------------------------
-- $Id: generic_ram-c.vhd,v 1.1 2005/12/17 02:11:40 arnim Exp $
-------------------------------------------------------------------------------

configuration generic_ram_rtl_c0 of generic_ram is

  for rtl
  end for;

end generic_ram_rtl_c0;
