
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity os_5200 is
port(
        clock:in std_logic;
        address:in std_logic_vector(10 downto 0);
        q:out std_logic_vector(7 downto 0)
);
end os_5200;

architecture syn of os_5200 is
        type rom_type is array(0 to 2047) of std_logic_vector(7 downto 0);
        signal ROM:rom_type:=
(
	X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"18",
X"18",
X"00",
X"18",
X"00",
X"00",
X"66",
X"66",
X"66",
X"00",
X"00",
X"00",
X"00",
X"00",
X"66",
X"ff",
X"66",
X"66",
X"ff",
X"66",
X"00",
X"18",
X"3e",
X"60",
X"3c",
X"06",
X"7c",
X"18",
X"00",
X"00",
X"66",
X"6c",
X"18",
X"30",
X"66",
X"46",
X"00",
X"1c",
X"36",
X"1c",
X"38",
X"6f",
X"66",
X"3b",
X"00",
X"00",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"00",
X"00",
X"0e",
X"1c",
X"18",
X"18",
X"1c",
X"0e",
X"00",
X"00",
X"70",
X"38",
X"18",
X"18",
X"38",
X"70",
X"00",
X"00",
X"66",
X"3c",
X"ff",
X"3c",
X"66",
X"00",
X"00",
X"00",
X"18",
X"18",
X"7e",
X"18",
X"18",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"30",
X"00",
X"00",
X"00",
X"7e",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"00",
X"00",
X"06",
X"0c",
X"18",
X"30",
X"60",
X"40",
X"00",
X"00",
X"3c",
X"66",
X"6e",
X"76",
X"66",
X"3c",
X"00",
X"00",
X"18",
X"38",
X"18",
X"18",
X"18",
X"7e",
X"00",
X"00",
X"3c",
X"66",
X"0c",
X"18",
X"30",
X"7e",
X"00",
X"00",
X"7e",
X"0c",
X"18",
X"0c",
X"66",
X"3c",
X"00",
X"00",
X"0c",
X"1c",
X"3c",
X"6c",
X"7e",
X"0c",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"06",
X"66",
X"3c",
X"00",
X"00",
X"3c",
X"60",
X"7c",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"7e",
X"06",
X"0c",
X"18",
X"30",
X"30",
X"00",
X"00",
X"3c",
X"66",
X"3c",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"3c",
X"66",
X"3e",
X"06",
X"0c",
X"38",
X"00",
X"00",
X"00",
X"18",
X"18",
X"00",
X"18",
X"18",
X"00",
X"00",
X"00",
X"18",
X"18",
X"00",
X"18",
X"18",
X"30",
X"06",
X"0c",
X"18",
X"30",
X"18",
X"0c",
X"06",
X"00",
X"00",
X"00",
X"7e",
X"00",
X"00",
X"7e",
X"00",
X"00",
X"60",
X"30",
X"18",
X"0c",
X"18",
X"30",
X"60",
X"00",
X"00",
X"3c",
X"66",
X"0c",
X"18",
X"00",
X"18",
X"00",
X"00",
X"3c",
X"66",
X"6e",
X"6e",
X"60",
X"3e",
X"00",
X"00",
X"18",
X"3c",
X"66",
X"66",
X"7e",
X"66",
X"00",
X"00",
X"7c",
X"66",
X"7c",
X"66",
X"66",
X"7c",
X"00",
X"00",
X"3c",
X"66",
X"60",
X"60",
X"66",
X"3c",
X"00",
X"00",
X"78",
X"6c",
X"66",
X"66",
X"6c",
X"78",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"60",
X"60",
X"7e",
X"00",
X"00",
X"7e",
X"60",
X"7c",
X"60",
X"60",
X"60",
X"00",
X"00",
X"3e",
X"60",
X"60",
X"6e",
X"66",
X"3e",
X"00",
X"00",
X"66",
X"66",
X"7e",
X"66",
X"66",
X"66",
X"00",
X"00",
X"7e",
X"18",
X"18",
X"18",
X"18",
X"7e",
X"00",
X"00",
X"06",
X"06",
X"06",
X"06",
X"66",
X"3c",
X"00",
X"00",
X"66",
X"6c",
X"78",
X"78",
X"6c",
X"66",
X"00",
X"00",
X"60",
X"60",
X"60",
X"60",
X"60",
X"7e",
X"00",
X"00",
X"63",
X"77",
X"7f",
X"6b",
X"63",
X"63",
X"00",
X"00",
X"66",
X"76",
X"7e",
X"7e",
X"6e",
X"66",
X"00",
X"00",
X"3c",
X"66",
X"66",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"7c",
X"60",
X"60",
X"00",
X"00",
X"3c",
X"66",
X"66",
X"66",
X"6c",
X"36",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"7c",
X"6c",
X"66",
X"00",
X"00",
X"3c",
X"60",
X"3c",
X"06",
X"06",
X"3c",
X"00",
X"00",
X"7e",
X"18",
X"18",
X"18",
X"18",
X"18",
X"00",
X"00",
X"66",
X"66",
X"66",
X"66",
X"66",
X"7e",
X"00",
X"00",
X"66",
X"66",
X"66",
X"66",
X"3c",
X"18",
X"00",
X"00",
X"63",
X"63",
X"6b",
X"7f",
X"77",
X"63",
X"00",
X"00",
X"66",
X"66",
X"3c",
X"3c",
X"66",
X"66",
X"00",
X"00",
X"66",
X"66",
X"3c",
X"18",
X"18",
X"18",
X"00",
X"00",
X"7e",
X"0c",
X"18",
X"30",
X"60",
X"7e",
X"00",
X"00",
X"1e",
X"18",
X"18",
X"18",
X"18",
X"1e",
X"00",
X"00",
X"40",
X"60",
X"30",
X"18",
X"0c",
X"06",
X"00",
X"00",
X"78",
X"18",
X"18",
X"18",
X"18",
X"78",
X"00",
X"00",
X"08",
X"1c",
X"36",
X"63",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"00",
X"00",
X"36",
X"7f",
X"7f",
X"3e",
X"1c",
X"08",
X"00",
X"18",
X"18",
X"18",
X"1f",
X"1f",
X"18",
X"18",
X"18",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"18",
X"18",
X"18",
X"f8",
X"f8",
X"00",
X"00",
X"00",
X"18",
X"18",
X"18",
X"f8",
X"f8",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"f8",
X"f8",
X"18",
X"18",
X"18",
X"03",
X"07",
X"0e",
X"1c",
X"38",
X"70",
X"e0",
X"c0",
X"c0",
X"e0",
X"70",
X"38",
X"1c",
X"0e",
X"07",
X"03",
X"01",
X"03",
X"07",
X"0f",
X"1f",
X"3f",
X"7f",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"0f",
X"0f",
X"0f",
X"0f",
X"80",
X"c0",
X"e0",
X"f0",
X"f8",
X"fc",
X"fe",
X"ff",
X"0f",
X"0f",
X"0f",
X"0f",
X"00",
X"00",
X"00",
X"00",
X"f0",
X"f0",
X"f0",
X"f0",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"f0",
X"f0",
X"f0",
X"f0",
X"00",
X"1c",
X"1c",
X"77",
X"77",
X"08",
X"1c",
X"00",
X"00",
X"00",
X"00",
X"1f",
X"1f",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"18",
X"18",
X"18",
X"ff",
X"ff",
X"18",
X"18",
X"18",
X"00",
X"00",
X"3c",
X"7e",
X"7e",
X"7e",
X"3c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"c0",
X"c0",
X"c0",
X"c0",
X"c0",
X"c0",
X"c0",
X"c0",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"18",
X"18",
X"18",
X"1f",
X"1f",
X"00",
X"00",
X"00",
X"78",
X"60",
X"78",
X"60",
X"7e",
X"18",
X"1e",
X"00",
X"00",
X"18",
X"3c",
X"7e",
X"18",
X"18",
X"18",
X"00",
X"00",
X"18",
X"18",
X"18",
X"7e",
X"3c",
X"18",
X"00",
X"00",
X"18",
X"30",
X"7e",
X"30",
X"18",
X"00",
X"00",
X"00",
X"18",
X"0c",
X"7e",
X"0c",
X"18",
X"00",
X"00",
X"00",
X"18",
X"3c",
X"7e",
X"7e",
X"3c",
X"18",
X"00",
X"00",
X"00",
X"3c",
X"06",
X"3e",
X"66",
X"3e",
X"00",
X"00",
X"60",
X"60",
X"7c",
X"66",
X"66",
X"7c",
X"00",
X"00",
X"00",
X"3c",
X"60",
X"60",
X"60",
X"3c",
X"00",
X"00",
X"06",
X"06",
X"3e",
X"66",
X"66",
X"3e",
X"00",
X"00",
X"00",
X"3c",
X"66",
X"7e",
X"60",
X"3c",
X"00",
X"00",
X"0e",
X"18",
X"3e",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"3e",
X"66",
X"66",
X"3e",
X"06",
X"7c",
X"00",
X"60",
X"60",
X"7c",
X"66",
X"66",
X"66",
X"00",
X"00",
X"18",
X"00",
X"38",
X"18",
X"18",
X"3c",
X"00",
X"00",
X"06",
X"00",
X"06",
X"06",
X"06",
X"06",
X"3c",
X"00",
X"60",
X"60",
X"6c",
X"78",
X"6c",
X"66",
X"00",
X"00",
X"38",
X"18",
X"18",
X"18",
X"18",
X"3c",
X"00",
X"00",
X"00",
X"66",
X"7f",
X"7f",
X"6b",
X"63",
X"00",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"66",
X"66",
X"00",
X"00",
X"00",
X"3c",
X"66",
X"66",
X"66",
X"3c",
X"00",
X"00",
X"00",
X"7c",
X"66",
X"66",
X"7c",
X"60",
X"60",
X"00",
X"00",
X"3e",
X"66",
X"66",
X"3e",
X"06",
X"06",
X"00",
X"00",
X"7c",
X"66",
X"60",
X"60",
X"60",
X"00",
X"00",
X"00",
X"3e",
X"60",
X"3c",
X"06",
X"7c",
X"00",
X"00",
X"18",
X"7e",
X"18",
X"18",
X"18",
X"0e",
X"00",
X"00",
X"00",
X"66",
X"66",
X"66",
X"66",
X"3e",
X"00",
X"00",
X"00",
X"66",
X"66",
X"66",
X"3c",
X"18",
X"00",
X"00",
X"00",
X"63",
X"6b",
X"7f",
X"3e",
X"36",
X"00",
X"00",
X"00",
X"66",
X"3c",
X"18",
X"3c",
X"66",
X"00",
X"00",
X"00",
X"66",
X"66",
X"66",
X"3e",
X"0c",
X"78",
X"00",
X"00",
X"7e",
X"0c",
X"18",
X"30",
X"7e",
X"00",
X"00",
X"18",
X"3c",
X"7e",
X"7e",
X"18",
X"3c",
X"00",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"00",
X"7e",
X"78",
X"7c",
X"6e",
X"66",
X"06",
X"00",
X"08",
X"18",
X"38",
X"78",
X"38",
X"18",
X"08",
X"00",
X"10",
X"18",
X"1c",
X"1e",
X"1c",
X"18",
X"10",
X"00",
X"6c",
X"00",
X"02",
X"48",
X"a9",
X"20",
X"2c",
X"0e",
X"e8",
X"d0",
X"0d",
X"a9",
X"df",
X"8d",
X"0e",
X"e8",
X"a5",
X"00",
X"8d",
X"0e",
X"e8",
X"6c",
X"10",
X"02",
X"10",
X"6e",
X"50",
X"79",
X"a9",
X"10",
X"2d",
X"0e",
X"e8",
X"d0",
X"0d",
X"a9",
X"ef",
X"8d",
X"0e",
X"e8",
X"a5",
X"00",
X"8d",
X"0e",
X"e8",
X"6c",
X"12",
X"02",
X"a9",
X"08",
X"25",
X"00",
X"f0",
X"12",
X"2d",
X"0e",
X"e8",
X"d0",
X"0d",
X"a9",
X"f7",
X"8d",
X"0e",
X"e8",
X"a5",
X"00",
X"8d",
X"0e",
X"e8",
X"6c",
X"14",
X"02",
X"ad",
X"0e",
X"e8",
X"6a",
X"b0",
X"0d",
X"a9",
X"fe",
X"8d",
X"0e",
X"e8",
X"a5",
X"00",
X"8d",
X"0e",
X"e8",
X"6c",
X"16",
X"02",
X"6a",
X"b0",
X"0d",
X"a9",
X"fd",
X"8d",
X"0e",
X"e8",
X"a5",
X"00",
X"8d",
X"0e",
X"e8",
X"6c",
X"18",
X"02",
X"6a",
X"b0",
X"0d",
X"a9",
X"fb",
X"8d",
X"0e",
X"e8",
X"a5",
X"00",
X"8d",
X"0e",
X"e8",
X"6c",
X"1a",
X"02",
X"8a",
X"48",
X"ba",
X"bd",
X"03",
X"01",
X"29",
X"10",
X"f0",
X"2f",
X"6c",
X"0e",
X"02",
X"a9",
X"7f",
X"8d",
X"0e",
X"e8",
X"a5",
X"00",
X"8d",
X"0e",
X"e8",
X"6c",
X"0c",
X"02",
X"a9",
X"bf",
X"8d",
X"0e",
X"e8",
X"a5",
X"00",
X"8d",
X"0e",
X"e8",
X"6c",
X"08",
X"02",
X"2c",
X"0f",
X"d4",
X"8d",
X"0f",
X"d4",
X"30",
X"05",
X"50",
X"0b",
X"6c",
X"02",
X"02",
X"6c",
X"06",
X"02",
X"68",
X"a8",
X"68",
X"aa",
X"68",
X"40",
X"48",
X"8a",
X"48",
X"98",
X"48",
X"e6",
X"02",
X"d0",
X"04",
X"e6",
X"04",
X"e6",
X"01",
X"a5",
X"03",
X"d0",
X"e9",
X"a5",
X"06",
X"8d",
X"03",
X"d4",
X"a5",
X"05",
X"8d",
X"02",
X"d4",
X"a5",
X"07",
X"8d",
X"00",
X"d4",
X"a4",
X"04",
X"10",
X"04",
X"a0",
X"80",
X"84",
X"04",
X"a2",
X"08",
X"b5",
X"08",
X"c0",
X"80",
X"90",
X"04",
X"45",
X"01",
X"29",
X"f6",
X"9d",
X"12",
X"c0",
X"ca",
X"10",
X"f0",
X"a2",
X"07",
X"bd",
X"00",
X"e8",
X"95",
X"11",
X"ca",
X"10",
X"f8",
X"8d",
X"0b",
X"e8",
X"6c",
X"04",
X"02",
X"8a",
X"48",
X"98",
X"48",
X"ad",
X"09",
X"e8",
X"4a",
X"29",
X"0f",
X"aa",
X"bd",
X"13",
X"fd",
X"6c",
X"0a",
X"02",
X"ff",
X"0b",
X"00",
X"0a",
X"0e",
X"09",
X"08",
X"07",
X"0d",
X"06",
X"05",
X"04",
X"0c",
X"03",
X"02",
X"01",
X"78",
X"d8",
X"a2",
X"ff",
X"9a",
X"ad",
X"fd",
X"bf",
X"c9",
X"ff",
X"d0",
X"03",
X"6c",
X"fe",
X"bf",
X"e8",
X"8a",
X"9d",
X"00",
X"e8",
X"9d",
X"00",
X"c0",
X"9d",
X"00",
X"d4",
X"95",
X"00",
X"e8",
X"d0",
X"f2",
X"a9",
X"f8",
X"8d",
X"09",
X"d4",
X"a2",
X"0b",
X"bd",
X"95",
X"fe",
X"9d",
X"00",
X"02",
X"ca",
X"10",
X"f7",
X"a9",
X"3c",
X"85",
X"12",
X"a9",
X"00",
X"85",
X"11",
X"a2",
X"0c",
X"a8",
X"91",
X"11",
X"88",
X"d0",
X"fb",
X"c6",
X"12",
X"ca",
X"10",
X"f6",
X"a9",
X"0d",
X"a2",
X"4d",
X"9d",
X"07",
X"20",
X"ca",
X"10",
X"fa",
X"a2",
X"06",
X"bd",
X"c8",
X"fe",
X"9d",
X"00",
X"20",
X"ca",
X"10",
X"f7",
X"a2",
X"04",
X"bd",
X"cf",
X"fe",
X"9d",
X"55",
X"20",
X"ca",
X"10",
X"f7",
X"a9",
X"00",
X"85",
X"05",
X"a9",
X"20",
X"85",
X"06",
X"a9",
X"22",
X"85",
X"07",
X"a9",
X"30",
X"a8",
X"a9",
X"28",
X"a2",
X"36",
X"9d",
X"00",
X"11",
X"48",
X"98",
X"9d",
X"00",
X"10",
X"68",
X"ca",
X"30",
X"08",
X"18",
X"69",
X"28",
X"90",
X"ef",
X"c8",
X"b0",
X"ec",
X"a2",
X"13",
X"86",
X"17",
X"e8",
X"86",
X"18",
X"a9",
X"20",
X"85",
X"13",
X"a9",
X"01",
X"85",
X"15",
X"a9",
X"40",
X"85",
X"16",
X"c6",
X"13",
X"30",
X"3e",
X"a6",
X"13",
X"bd",
X"e8",
X"fe",
X"85",
X"14",
X"bd",
X"08",
X"ff",
X"aa",
X"e4",
X"14",
X"f0",
X"1d",
X"bd",
X"00",
X"11",
X"85",
X"11",
X"bd",
X"00",
X"10",
X"85",
X"12",
X"a4",
X"17",
X"a5",
X"15",
X"11",
X"11",
X"91",
X"11",
X"a4",
X"18",
X"a5",
X"16",
X"11",
X"11",
X"91",
X"11",
X"e8",
X"d0",
X"df",
X"06",
X"15",
X"06",
X"15",
X"b0",
X"06",
X"46",
X"16",
X"46",
X"16",
X"90",
X"c4",
X"c6",
X"17",
X"e6",
X"18",
X"b0",
X"b6",
X"a9",
X"11",
X"85",
X"11",
X"a9",
X"39",
X"85",
X"12",
X"a9",
X"13",
X"85",
X"13",
X"a9",
X"00",
X"85",
X"15",
X"a9",
X"01",
X"a0",
X"0a",
X"85",
X"18",
X"a6",
X"15",
X"e6",
X"15",
X"bd",
X"28",
X"ff",
X"f0",
X"2a",
X"aa",
X"29",
X"0f",
X"85",
X"16",
X"8a",
X"4a",
X"4a",
X"4a",
X"4a",
X"aa",
X"a5",
X"18",
X"0a",
X"0a",
X"90",
X"05",
X"91",
X"11",
X"c8",
X"a9",
X"01",
X"ca",
X"10",
X"f4",
X"a6",
X"16",
X"38",
X"2a",
X"0a",
X"90",
X"05",
X"91",
X"11",
X"c8",
X"a9",
X"01",
X"ca",
X"10",
X"f3",
X"30",
X"cb",
X"a5",
X"18",
X"0a",
X"0a",
X"90",
X"fc",
X"91",
X"11",
X"a5",
X"11",
X"18",
X"69",
X"28",
X"85",
X"11",
X"90",
X"02",
X"e6",
X"12",
X"c6",
X"13",
X"10",
X"b0",
X"a2",
X"13",
X"bd",
X"d4",
X"fe",
X"9d",
X"94",
X"3c",
X"bd",
X"e8",
X"bf",
X"9d",
X"80",
X"3c",
X"ca",
X"10",
X"f1",
X"ad",
X"fc",
X"bf",
X"8d",
X"a0",
X"3c",
X"ad",
X"fd",
X"bf",
X"8d",
X"a1",
X"3c",
X"a9",
X"0f",
X"85",
X"0d",
X"a9",
X"c0",
X"8d",
X"0e",
X"d4",
X"a9",
X"02",
X"8d",
X"0f",
X"e8",
X"e4",
X"02",
X"d0",
X"fc",
X"6c",
X"fe",
X"bf",
X"03",
X"fc",
X"b8",
X"fc",
X"b2",
X"fc",
X"a1",
X"fe",
X"02",
X"fd",
X"b2",
X"fc",
X"48",
X"8a",
X"48",
X"98",
X"48",
X"a6",
X"08",
X"a0",
X"72",
X"e0",
X"10",
X"b0",
X"02",
X"a2",
X"fe",
X"8e",
X"0a",
X"d4",
X"8e",
X"16",
X"c0",
X"ca",
X"ca",
X"88",
X"d0",
X"ef",
X"e6",
X"08",
X"a0",
X"10",
X"c4",
X"08",
X"90",
X"02",
X"84",
X"08",
X"4c",
X"b2",
X"fc",
X"70",
X"70",
X"70",
X"4d",
X"00",
X"30",
X"8d",
X"07",
X"07",
X"41",
X"00",
X"20",
X"63",
X"6f",
X"70",
X"79",
X"72",
X"69",
X"67",
X"68",
X"74",
X"00",
X"51",
X"59",
X"58",
X"51",
X"00",
X"61",
X"74",
X"61",
X"72",
X"69",
X"08",
X"08",
X"08",
X"09",
X"09",
X"09",
X"0a",
X"0a",
X"0b",
X"0b",
X"0c",
X"0d",
X"0e",
X"0f",
X"10",
X"11",
X"12",
X"14",
X"16",
X"19",
X"1c",
X"1f",
X"36",
X"36",
X"36",
X"36",
X"00",
X"00",
X"36",
X"36",
X"36",
X"36",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"02",
X"02",
X"03",
X"03",
X"04",
X"05",
X"06",
X"07",
X"08",
X"09",
X"0a",
X"0b",
X"0c",
X"0e",
X"10",
X"13",
X"16",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"92",
X"4e",
X"42",
X"97",
X"52",
X"00",
X"84",
X"3e",
X"34",
X"79",
X"42",
X"00",
X"76",
X"2e",
X"26",
X"5b",
X"32",
X"00",
X"76",
X"82",
X"86",
X"53",
X"43",
X"22",
X"00",
X"63",
X"03",
X"72",
X"73",
X"03",
X"42",
X"63",
X"12",
X"00",
X"62",
X"22",
X"72",
X"72",
X"22",
X"42",
X"72",
X"12",
X"00",
X"62",
X"22",
X"72",
X"72",
X"22",
X"42",
X"72",
X"12",
X"00",
X"52",
X"42",
X"62",
X"62",
X"42",
X"32",
X"62",
X"22",
X"00",
X"52",
X"42",
X"62",
X"62",
X"42",
X"32",
X"52",
X"32",
X"00",
X"52",
X"42",
X"62",
X"62",
X"42",
X"32",
X"06",
X"42",
X"00",
X"43",
X"43",
X"52",
X"53",
X"43",
X"22",
X"05",
X"52",
X"00",
X"42",
X"62",
X"52",
X"52",
X"62",
X"22",
X"05",
X"52",
X"00",
X"42",
X"62",
X"52",
X"52",
X"62",
X"22",
X"42",
X"42",
X"00",
X"3e",
X"42",
X"4e",
X"12",
X"42",
X"42",
X"00",
X"3e",
X"42",
X"4e",
X"12",
X"52",
X"32",
X"00",
X"3e",
X"42",
X"4e",
X"12",
X"52",
X"32",
X"00",
X"23",
X"83",
X"32",
X"33",
X"83",
X"02",
X"62",
X"22",
X"00",
X"22",
X"a2",
X"32",
X"32",
X"a2",
X"02",
X"62",
X"22",
X"00",
X"22",
X"a2",
X"32",
X"32",
X"a2",
X"02",
X"72",
X"12",
X"00",
X"22",
X"a2",
X"32",
X"32",
X"a2",
X"02",
X"72",
X"12",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"52",
X"4a",
X"5a",
X"20",
X"31",
X"39",
X"38",
X"32",
X"00",
X"a2",
X"fc",
X"23",
X"fd",
X"00",
X"fc"

);
        signal rdata:std_logic_vector(7 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
