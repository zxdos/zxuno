
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity os2 is
port(
        clock:in std_logic;
        address:in std_logic_vector(10 downto 0);
        q:out std_logic_vector(7 downto 0)
);
end os2;

architecture syn of os2 is
        type rom_type is array(0 to 2047) of std_logic_vector(7 downto 0);
        signal ROM:rom_type:=
(
	X"20",
X"a1",
X"db",
X"20",
X"bb",
X"db",
X"b0",
X"39",
X"a2",
X"ed",
X"a0",
X"04",
X"20",
X"48",
X"da",
X"a2",
X"ff",
X"86",
X"f1",
X"20",
X"44",
X"da",
X"f0",
X"04",
X"a9",
X"ff",
X"85",
X"f0",
X"20",
X"94",
X"db",
X"b0",
X"21",
X"48",
X"a6",
X"d5",
X"d0",
X"11",
X"20",
X"eb",
X"db",
X"68",
X"05",
X"d9",
X"85",
X"d9",
X"a6",
X"f1",
X"30",
X"e6",
X"e8",
X"86",
X"f1",
X"d0",
X"e1",
X"68",
X"a6",
X"f1",
X"10",
X"02",
X"e6",
X"ed",
X"4c",
X"18",
X"d8",
X"60",
X"c9",
X"2e",
X"f0",
X"14",
X"c9",
X"45",
X"f0",
X"19",
X"a6",
X"f0",
X"d0",
X"68",
X"c9",
X"2b",
X"f0",
X"c6",
X"c9",
X"2d",
X"f0",
X"00",
X"85",
X"ee",
X"f0",
X"be",
X"a6",
X"f1",
X"10",
X"58",
X"e8",
X"86",
X"f1",
X"f0",
X"b5",
X"a5",
X"f2",
X"85",
X"ec",
X"20",
X"94",
X"db",
X"b0",
X"37",
X"aa",
X"a5",
X"ed",
X"48",
X"86",
X"ed",
X"20",
X"94",
X"db",
X"b0",
X"17",
X"48",
X"a5",
X"ed",
X"0a",
X"85",
X"ed",
X"0a",
X"0a",
X"65",
X"ed",
X"85",
X"ed",
X"68",
X"18",
X"65",
X"ed",
X"85",
X"ed",
X"a4",
X"f2",
X"20",
X"9d",
X"db",
X"a5",
X"ef",
X"f0",
X"09",
X"a5",
X"ed",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"85",
X"ed",
X"68",
X"18",
X"65",
X"ed",
X"85",
X"ed",
X"d0",
X"13",
X"c9",
X"2b",
X"f0",
X"06",
X"c9",
X"2d",
X"d0",
X"07",
X"85",
X"ef",
X"20",
X"94",
X"db",
X"90",
X"ba",
X"a5",
X"ec",
X"85",
X"f2",
X"c6",
X"f2",
X"a5",
X"ed",
X"a6",
X"f1",
X"30",
X"05",
X"f0",
X"03",
X"38",
X"e5",
X"f1",
X"48",
X"2a",
X"68",
X"6a",
X"85",
X"ed",
X"90",
X"03",
X"20",
X"eb",
X"db",
X"a5",
X"ed",
X"18",
X"69",
X"44",
X"85",
X"d4",
X"20",
X"00",
X"dc",
X"b0",
X"0b",
X"a6",
X"ee",
X"f0",
X"06",
X"a5",
X"d4",
X"09",
X"80",
X"85",
X"d4",
X"18",
X"60",
X"20",
X"51",
X"da",
X"a9",
X"30",
X"8d",
X"7f",
X"05",
X"a5",
X"d4",
X"f0",
X"28",
X"29",
X"7f",
X"c9",
X"3f",
X"90",
X"28",
X"c9",
X"45",
X"b0",
X"24",
X"38",
X"e9",
X"3f",
X"20",
X"70",
X"dc",
X"20",
X"a4",
X"dc",
X"09",
X"80",
X"9d",
X"80",
X"05",
X"ad",
X"80",
X"05",
X"c9",
X"2e",
X"f0",
X"03",
X"4c",
X"88",
X"d9",
X"20",
X"c1",
X"dc",
X"4c",
X"9c",
X"d9",
X"a9",
X"b0",
X"8d",
X"80",
X"05",
X"60",
X"a9",
X"01",
X"20",
X"70",
X"dc",
X"20",
X"a4",
X"dc",
X"e8",
X"86",
X"f2",
X"a5",
X"d4",
X"0a",
X"38",
X"e9",
X"80",
X"ae",
X"80",
X"05",
X"e0",
X"30",
X"f0",
X"17",
X"ae",
X"81",
X"05",
X"ac",
X"82",
X"05",
X"8e",
X"82",
X"05",
X"8c",
X"81",
X"05",
X"a6",
X"f2",
X"e0",
X"02",
X"d0",
X"02",
X"e6",
X"f2",
X"18",
X"69",
X"01",
X"85",
X"ed",
X"a9",
X"45",
X"a4",
X"f2",
X"20",
X"9f",
X"dc",
X"84",
X"f2",
X"a5",
X"ed",
X"10",
X"0b",
X"a9",
X"00",
X"38",
X"e5",
X"ed",
X"85",
X"ed",
X"a9",
X"2d",
X"d0",
X"02",
X"a9",
X"2b",
X"20",
X"9f",
X"dc",
X"a2",
X"00",
X"a5",
X"ed",
X"38",
X"e9",
X"0a",
X"90",
X"03",
X"e8",
X"d0",
X"f8",
X"18",
X"69",
X"0a",
X"48",
X"8a",
X"20",
X"9d",
X"dc",
X"68",
X"09",
X"80",
X"20",
X"9d",
X"dc",
X"ad",
X"80",
X"05",
X"c9",
X"30",
X"d0",
X"0d",
X"18",
X"a5",
X"f3",
X"69",
X"01",
X"85",
X"f3",
X"a5",
X"f4",
X"69",
X"00",
X"85",
X"f4",
X"a5",
X"d4",
X"10",
X"09",
X"20",
X"c1",
X"dc",
X"a0",
X"00",
X"a9",
X"2d",
X"91",
X"f3",
X"60",
X"a5",
X"d4",
X"85",
X"f8",
X"a5",
X"d5",
X"85",
X"f7",
X"20",
X"44",
X"da",
X"f8",
X"a0",
X"10",
X"06",
X"f8",
X"26",
X"f7",
X"a2",
X"03",
X"b5",
X"d4",
X"75",
X"d4",
X"95",
X"d4",
X"ca",
X"d0",
X"f7",
X"88",
X"d0",
X"ee",
X"d8",
X"a9",
X"42",
X"85",
X"d4",
X"4c",
X"00",
X"dc",
X"a9",
X"00",
X"85",
X"f7",
X"85",
X"f8",
X"a5",
X"d4",
X"30",
X"66",
X"c9",
X"43",
X"b0",
X"62",
X"38",
X"e9",
X"40",
X"90",
X"3f",
X"69",
X"00",
X"0a",
X"85",
X"f5",
X"20",
X"5a",
X"da",
X"b0",
X"53",
X"a5",
X"f7",
X"85",
X"f9",
X"a5",
X"f8",
X"85",
X"fa",
X"20",
X"5a",
X"da",
X"b0",
X"46",
X"20",
X"5a",
X"da",
X"b0",
X"41",
X"18",
X"a5",
X"f8",
X"65",
X"fa",
X"85",
X"f8",
X"a5",
X"f7",
X"65",
X"f9",
X"85",
X"f7",
X"b0",
X"32",
X"20",
X"b9",
X"dc",
X"18",
X"65",
X"f8",
X"85",
X"f8",
X"a5",
X"f7",
X"69",
X"00",
X"b0",
X"24",
X"85",
X"f7",
X"c6",
X"f5",
X"d0",
X"c6",
X"20",
X"b9",
X"dc",
X"c9",
X"05",
X"90",
X"0d",
X"18",
X"a5",
X"f8",
X"69",
X"01",
X"85",
X"f8",
X"a5",
X"f7",
X"69",
X"00",
X"85",
X"f7",
X"a5",
X"f8",
X"85",
X"d4",
X"a5",
X"f7",
X"85",
X"d5",
X"18",
X"60",
X"38",
X"60",
X"a2",
X"d4",
X"a0",
X"06",
X"a9",
X"00",
X"95",
X"00",
X"e8",
X"88",
X"d0",
X"fa",
X"60",
X"a9",
X"05",
X"85",
X"f4",
X"a9",
X"80",
X"85",
X"f3",
X"60",
X"18",
X"26",
X"f8",
X"26",
X"f7",
X"60",
X"a5",
X"e0",
X"49",
X"80",
X"85",
X"e0",
X"a5",
X"e0",
X"29",
X"7f",
X"85",
X"f7",
X"a5",
X"d4",
X"29",
X"7f",
X"38",
X"e5",
X"f7",
X"10",
X"10",
X"a2",
X"05",
X"b5",
X"d4",
X"b4",
X"e0",
X"95",
X"e0",
X"98",
X"95",
X"d4",
X"ca",
X"10",
X"f4",
X"30",
X"e1",
X"f0",
X"07",
X"c9",
X"05",
X"b0",
X"19",
X"20",
X"3e",
X"dc",
X"f8",
X"a5",
X"d4",
X"45",
X"e0",
X"30",
X"1e",
X"a2",
X"04",
X"18",
X"b5",
X"d5",
X"75",
X"e1",
X"95",
X"d5",
X"ca",
X"10",
X"f7",
X"d8",
X"b0",
X"03",
X"4c",
X"00",
X"dc",
X"a9",
X"01",
X"20",
X"3a",
X"dc",
X"a9",
X"01",
X"85",
X"d5",
X"4c",
X"00",
X"dc",
X"a2",
X"04",
X"38",
X"b5",
X"d5",
X"f5",
X"e1",
X"95",
X"d5",
X"ca",
X"10",
X"f7",
X"90",
X"04",
X"d8",
X"4c",
X"00",
X"dc",
X"a5",
X"d4",
X"49",
X"80",
X"85",
X"d4",
X"38",
X"a2",
X"04",
X"a9",
X"00",
X"f5",
X"d5",
X"95",
X"d5",
X"ca",
X"10",
X"f7",
X"d8",
X"4c",
X"00",
X"dc",
X"a5",
X"d4",
X"f0",
X"45",
X"a5",
X"e0",
X"f0",
X"3e",
X"20",
X"cf",
X"dc",
X"38",
X"e9",
X"40",
X"38",
X"65",
X"e0",
X"30",
X"38",
X"20",
X"e0",
X"dc",
X"a5",
X"df",
X"29",
X"0f",
X"85",
X"f6",
X"c6",
X"f6",
X"30",
X"06",
X"20",
X"01",
X"dd",
X"4c",
X"f7",
X"da",
X"a5",
X"df",
X"4a",
X"4a",
X"4a",
X"4a",
X"85",
X"f6",
X"c6",
X"f6",
X"30",
X"06",
X"20",
X"05",
X"dd",
X"4c",
X"09",
X"db",
X"20",
X"62",
X"dc",
X"c6",
X"f5",
X"d0",
X"d7",
X"a5",
X"ed",
X"85",
X"d4",
X"4c",
X"04",
X"dc",
X"20",
X"44",
X"da",
X"18",
X"60",
X"38",
X"60",
X"a5",
X"e0",
X"f0",
X"fa",
X"a5",
X"d4",
X"f0",
X"f4",
X"20",
X"cf",
X"dc",
X"38",
X"e5",
X"e0",
X"18",
X"69",
X"40",
X"30",
X"eb",
X"20",
X"e0",
X"dc",
X"e6",
X"f5",
X"4c",
X"4e",
X"db",
X"a2",
X"00",
X"b5",
X"d5",
X"95",
X"d4",
X"e8",
X"e0",
X"0c",
X"d0",
X"f7",
X"a0",
X"05",
X"38",
X"f8",
X"b9",
X"da",
X"00",
X"f9",
X"e6",
X"00",
X"99",
X"da",
X"00",
X"88",
X"10",
X"f4",
X"d8",
X"90",
X"04",
X"e6",
X"d9",
X"d0",
X"e9",
X"20",
X"0f",
X"dd",
X"06",
X"d9",
X"06",
X"d9",
X"06",
X"d9",
X"06",
X"d9",
X"a0",
X"05",
X"38",
X"f8",
X"b9",
X"da",
X"00",
X"f9",
X"e0",
X"00",
X"99",
X"da",
X"00",
X"88",
X"10",
X"f4",
X"d8",
X"90",
X"04",
X"e6",
X"d9",
X"d0",
X"e9",
X"20",
X"09",
X"dd",
X"c6",
X"f5",
X"d0",
X"b5",
X"20",
X"62",
X"dc",
X"4c",
X"1a",
X"db",
X"20",
X"af",
X"db",
X"a4",
X"f2",
X"90",
X"02",
X"b1",
X"f3",
X"c8",
X"84",
X"f2",
X"60",
X"a4",
X"f2",
X"a9",
X"20",
X"d1",
X"f3",
X"d0",
X"03",
X"c8",
X"d0",
X"f9",
X"84",
X"f2",
X"60",
X"a4",
X"f2",
X"b1",
X"f3",
X"38",
X"e9",
X"30",
X"90",
X"18",
X"c9",
X"0a",
X"60",
X"a5",
X"f2",
X"48",
X"20",
X"94",
X"db",
X"90",
X"1f",
X"c9",
X"2e",
X"f0",
X"14",
X"c9",
X"2b",
X"f0",
X"07",
X"c9",
X"2d",
X"f0",
X"03",
X"68",
X"38",
X"60",
X"20",
X"94",
X"db",
X"90",
X"0b",
X"c9",
X"2e",
X"d0",
X"f4",
X"20",
X"94",
X"db",
X"90",
X"02",
X"b0",
X"ed",
X"68",
X"85",
X"f2",
X"18",
X"60",
X"a2",
X"e7",
X"d0",
X"02",
X"a2",
X"d5",
X"a0",
X"04",
X"18",
X"36",
X"04",
X"36",
X"03",
X"36",
X"02",
X"36",
X"01",
X"36",
X"00",
X"26",
X"ec",
X"88",
X"d0",
X"f0",
X"60",
X"a2",
X"00",
X"86",
X"da",
X"a2",
X"04",
X"a5",
X"d4",
X"f0",
X"2e",
X"a5",
X"d5",
X"d0",
X"1a",
X"a0",
X"00",
X"b9",
X"d6",
X"00",
X"99",
X"d5",
X"00",
X"c8",
X"c0",
X"05",
X"90",
X"f5",
X"c6",
X"d4",
X"ca",
X"d0",
X"ea",
X"a5",
X"d5",
X"d0",
X"04",
X"85",
X"d4",
X"18",
X"60",
X"a5",
X"d4",
X"29",
X"7f",
X"c9",
X"71",
X"90",
X"01",
X"60",
X"c9",
X"0f",
X"b0",
X"03",
X"20",
X"44",
X"da",
X"18",
X"60",
X"a2",
X"d4",
X"d0",
X"02",
X"a2",
X"e0",
X"86",
X"f9",
X"85",
X"f7",
X"85",
X"f8",
X"a0",
X"04",
X"b5",
X"04",
X"95",
X"05",
X"ca",
X"88",
X"d0",
X"f8",
X"a9",
X"00",
X"95",
X"05",
X"a6",
X"f9",
X"c6",
X"f7",
X"d0",
X"ec",
X"b5",
X"00",
X"18",
X"65",
X"f8",
X"95",
X"00",
X"60",
X"a2",
X"0a",
X"b5",
X"d4",
X"95",
X"d5",
X"ca",
X"10",
X"f9",
X"a9",
X"00",
X"85",
X"d4",
X"60",
X"85",
X"f7",
X"a2",
X"00",
X"a0",
X"00",
X"20",
X"93",
X"dc",
X"38",
X"e9",
X"01",
X"85",
X"f7",
X"b5",
X"d5",
X"4a",
X"4a",
X"4a",
X"4a",
X"20",
X"9d",
X"dc",
X"b5",
X"d5",
X"29",
X"0f",
X"20",
X"9d",
X"dc",
X"e8",
X"e0",
X"05",
X"90",
X"e3",
X"a5",
X"f7",
X"d0",
X"05",
X"a9",
X"2e",
X"20",
X"9f",
X"dc",
X"60",
X"09",
X"30",
X"99",
X"80",
X"05",
X"c8",
X"60",
X"a2",
X"0a",
X"bd",
X"80",
X"05",
X"c9",
X"2e",
X"f0",
X"07",
X"c9",
X"30",
X"d0",
X"07",
X"ca",
X"d0",
X"f2",
X"ca",
X"bd",
X"80",
X"05",
X"60",
X"20",
X"eb",
X"db",
X"a5",
X"ec",
X"29",
X"0f",
X"60",
X"38",
X"a5",
X"f3",
X"e9",
X"01",
X"85",
X"f3",
X"a5",
X"f4",
X"e9",
X"00",
X"85",
X"f4",
X"60",
X"a5",
X"d4",
X"45",
X"e0",
X"29",
X"80",
X"85",
X"ee",
X"06",
X"e0",
X"46",
X"e0",
X"a5",
X"d4",
X"29",
X"7f",
X"60",
X"05",
X"ee",
X"85",
X"ed",
X"a9",
X"00",
X"85",
X"d4",
X"85",
X"e0",
X"20",
X"28",
X"dd",
X"20",
X"e7",
X"db",
X"a5",
X"ec",
X"29",
X"0f",
X"85",
X"e6",
X"a9",
X"05",
X"85",
X"f5",
X"20",
X"34",
X"dd",
X"20",
X"44",
X"da",
X"60",
X"a2",
X"d9",
X"d0",
X"06",
X"a2",
X"d9",
X"d0",
X"08",
X"a2",
X"df",
X"a0",
X"e5",
X"d0",
X"04",
X"a2",
X"df",
X"a0",
X"eb",
X"a9",
X"05",
X"85",
X"f7",
X"18",
X"f8",
X"b5",
X"00",
X"79",
X"00",
X"00",
X"95",
X"00",
X"ca",
X"88",
X"c6",
X"f7",
X"10",
X"f3",
X"d8",
X"60",
X"a0",
X"05",
X"b9",
X"e0",
X"00",
X"99",
X"e6",
X"00",
X"88",
X"10",
X"f7",
X"60",
X"a0",
X"05",
X"b9",
X"d4",
X"00",
X"99",
X"da",
X"00",
X"88",
X"10",
X"f7",
X"60",
X"86",
X"fe",
X"84",
X"ff",
X"85",
X"ef",
X"a2",
X"e0",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"20",
X"b6",
X"dd",
X"a6",
X"fe",
X"a4",
X"ff",
X"20",
X"89",
X"dd",
X"c6",
X"ef",
X"f0",
X"2d",
X"20",
X"db",
X"da",
X"b0",
X"28",
X"18",
X"a5",
X"fe",
X"69",
X"06",
X"85",
X"fe",
X"90",
X"06",
X"a5",
X"ff",
X"69",
X"00",
X"85",
X"ff",
X"a6",
X"fe",
X"a4",
X"ff",
X"20",
X"98",
X"dd",
X"20",
X"66",
X"da",
X"b0",
X"0d",
X"c6",
X"ef",
X"f0",
X"09",
X"a2",
X"e0",
X"a0",
X"05",
X"20",
X"98",
X"dd",
X"30",
X"d3",
X"60",
X"86",
X"fc",
X"84",
X"fd",
X"a0",
X"05",
X"b1",
X"fc",
X"99",
X"d4",
X"00",
X"88",
X"10",
X"f8",
X"60",
X"86",
X"fc",
X"84",
X"fd",
X"a0",
X"05",
X"b1",
X"fc",
X"99",
X"e0",
X"00",
X"88",
X"10",
X"f8",
X"60",
X"86",
X"fc",
X"84",
X"fd",
X"a0",
X"05",
X"b9",
X"d4",
X"00",
X"91",
X"fc",
X"88",
X"10",
X"f8",
X"60",
X"a2",
X"05",
X"b5",
X"d4",
X"95",
X"e0",
X"ca",
X"10",
X"f9",
X"60",
X"a2",
X"89",
X"a0",
X"de",
X"20",
X"98",
X"dd",
X"20",
X"db",
X"da",
X"b0",
X"7f",
X"a9",
X"00",
X"85",
X"f1",
X"a5",
X"d4",
X"85",
X"f0",
X"29",
X"7f",
X"85",
X"d4",
X"38",
X"e9",
X"40",
X"30",
X"26",
X"c9",
X"04",
X"10",
X"6a",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"20",
X"d2",
X"d9",
X"a5",
X"d4",
X"85",
X"f1",
X"a5",
X"d5",
X"d0",
X"58",
X"20",
X"aa",
X"d9",
X"20",
X"b6",
X"dd",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"89",
X"dd",
X"20",
X"60",
X"da",
X"a9",
X"0a",
X"a2",
X"4d",
X"a0",
X"de",
X"20",
X"40",
X"dd",
X"20",
X"b6",
X"dd",
X"20",
X"db",
X"da",
X"a5",
X"f1",
X"f0",
X"23",
X"18",
X"6a",
X"85",
X"e0",
X"a9",
X"01",
X"90",
X"02",
X"a9",
X"10",
X"85",
X"e1",
X"a2",
X"04",
X"a9",
X"00",
X"95",
X"e2",
X"ca",
X"10",
X"fb",
X"a5",
X"e0",
X"18",
X"69",
X"40",
X"b0",
X"19",
X"30",
X"17",
X"85",
X"e0",
X"20",
X"db",
X"da",
X"a5",
X"f0",
X"10",
X"0d",
X"20",
X"b6",
X"dd",
X"a2",
X"8f",
X"a0",
X"de",
X"20",
X"89",
X"dd",
X"20",
X"28",
X"db",
X"60",
X"38",
X"60",
X"3d",
X"17",
X"94",
X"19",
X"00",
X"00",
X"3d",
X"57",
X"33",
X"05",
X"00",
X"00",
X"3e",
X"05",
X"54",
X"76",
X"62",
X"00",
X"3e",
X"32",
X"19",
X"62",
X"27",
X"00",
X"3f",
X"01",
X"68",
X"60",
X"30",
X"36",
X"3f",
X"07",
X"32",
X"03",
X"27",
X"41",
X"3f",
X"25",
X"43",
X"34",
X"56",
X"75",
X"3f",
X"66",
X"27",
X"37",
X"30",
X"50",
X"40",
X"01",
X"15",
X"12",
X"92",
X"55",
X"3f",
X"99",
X"99",
X"99",
X"99",
X"99",
X"3f",
X"43",
X"42",
X"94",
X"48",
X"19",
X"40",
X"01",
X"00",
X"00",
X"00",
X"00",
X"86",
X"fe",
X"84",
X"ff",
X"a2",
X"e0",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"a6",
X"fe",
X"a4",
X"ff",
X"20",
X"98",
X"dd",
X"20",
X"66",
X"da",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"a2",
X"e0",
X"a0",
X"05",
X"20",
X"89",
X"dd",
X"a6",
X"fe",
X"a4",
X"ff",
X"20",
X"98",
X"dd",
X"20",
X"60",
X"da",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"98",
X"dd",
X"20",
X"28",
X"db",
X"60",
X"a9",
X"01",
X"d0",
X"02",
X"a9",
X"00",
X"85",
X"f0",
X"a5",
X"d4",
X"10",
X"02",
X"38",
X"60",
X"a5",
X"d4",
X"85",
X"e0",
X"38",
X"e9",
X"40",
X"0a",
X"85",
X"f1",
X"a5",
X"d5",
X"29",
X"f0",
X"d0",
X"04",
X"a9",
X"01",
X"d0",
X"04",
X"e6",
X"f1",
X"a9",
X"10",
X"85",
X"e1",
X"a2",
X"04",
X"a9",
X"00",
X"95",
X"e2",
X"ca",
X"10",
X"fb",
X"20",
X"28",
X"db",
X"a2",
X"66",
X"a0",
X"df",
X"20",
X"95",
X"de",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"a7",
X"dd",
X"20",
X"b6",
X"dd",
X"20",
X"db",
X"da",
X"a9",
X"0a",
X"a2",
X"72",
X"a0",
X"df",
X"20",
X"40",
X"dd",
X"a2",
X"e6",
X"a0",
X"05",
X"20",
X"98",
X"dd",
X"20",
X"db",
X"da",
X"a2",
X"6c",
X"a0",
X"df",
X"20",
X"98",
X"dd",
X"20",
X"66",
X"da",
X"20",
X"b6",
X"dd",
X"a9",
X"00",
X"85",
X"d5",
X"a5",
X"f1",
X"85",
X"d4",
X"10",
X"07",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"85",
X"d4",
X"20",
X"aa",
X"d9",
X"24",
X"f1",
X"10",
X"06",
X"a9",
X"80",
X"05",
X"d4",
X"85",
X"d4",
X"20",
X"66",
X"da",
X"a5",
X"f0",
X"f0",
X"0a",
X"a2",
X"89",
X"a0",
X"de",
X"20",
X"98",
X"dd",
X"20",
X"28",
X"db",
X"18",
X"60",
X"40",
X"03",
X"16",
X"22",
X"77",
X"66",
X"3f",
X"50",
X"00",
X"00",
X"00",
X"00",
X"3f",
X"49",
X"15",
X"57",
X"11",
X"08",
X"bf",
X"51",
X"70",
X"49",
X"47",
X"08",
X"3f",
X"39",
X"20",
X"57",
X"61",
X"95",
X"bf",
X"04",
X"39",
X"63",
X"03",
X"55",
X"3f",
X"10",
X"09",
X"30",
X"12",
X"64",
X"3f",
X"09",
X"39",
X"08",
X"04",
X"60",
X"3f",
X"12",
X"42",
X"58",
X"47",
X"42",
X"3f",
X"17",
X"37",
X"12",
X"06",
X"08",
X"3f",
X"28",
X"95",
X"29",
X"71",
X"17",
X"3f",
X"86",
X"85",
X"88",
X"96",
X"44",
X"3e",
X"16",
X"05",
X"44",
X"49",
X"00",
X"be",
X"95",
X"68",
X"38",
X"45",
X"00",
X"3f",
X"02",
X"68",
X"79",
X"94",
X"16",
X"bf",
X"04",
X"92",
X"78",
X"90",
X"80",
X"3f",
X"07",
X"03",
X"15",
X"20",
X"00",
X"bf",
X"08",
X"92",
X"29",
X"12",
X"44",
X"3f",
X"11",
X"08",
X"40",
X"09",
X"11",
X"bf",
X"14",
X"28",
X"31",
X"56",
X"04",
X"3f",
X"19",
X"99",
X"98",
X"77",
X"44",
X"bf",
X"33",
X"33",
X"33",
X"31",
X"13",
X"3f",
X"99",
X"99",
X"99",
X"99",
X"99",
X"3f",
X"78",
X"53",
X"98",
X"16",
X"34",
X"98",
X"16",
X"34",
X"fc",
X"e0",
X"32",
X"50",
X"d9",
X"68",
X"11"

);
        signal rdata:std_logic_vector(7 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
