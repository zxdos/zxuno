-------------------------------------------------------------------------------
--
-- FPGA Colecovision
--
-- $Id: cv_addr_dec-c.vhd,v 1.2 2006/01/05 22:25:25 arnim Exp $
--
-------------------------------------------------------------------------------

configuration cv_addr_dec_rtl_c0 of cv_addr_dec is

  for rtl
  end for;

end cv_addr_dec_rtl_c0;
