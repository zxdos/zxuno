-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80d6",
     9 => x"c4080b0b",
    10 => x"80d6c808",
    11 => x"0b0b80d6",
    12 => x"cc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"d6cc0c0b",
    16 => x"0b80d6c8",
    17 => x"0c0b0b80",
    18 => x"d6c40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80d0ac",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80d6c470",
    57 => x"80e0fc27",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51a3cc",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80d6",
    65 => x"d40c9f0b",
    66 => x"80d6d80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"d6d808ff",
    70 => x"0580d6d8",
    71 => x"0c80d6d8",
    72 => x"088025e8",
    73 => x"3880d6d4",
    74 => x"08ff0580",
    75 => x"d6d40c80",
    76 => x"d6d40880",
    77 => x"25d03880",
    78 => x"0b80d6d8",
    79 => x"0c800b80",
    80 => x"d6d40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80d6d408",
   100 => x"25913882",
   101 => x"c82d80d6",
   102 => x"d408ff05",
   103 => x"80d6d40c",
   104 => x"838a0480",
   105 => x"d6d40880",
   106 => x"d6d80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80d6d408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"d6d80881",
   116 => x"0580d6d8",
   117 => x"0c80d6d8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80d6d8",
   121 => x"0c80d6d4",
   122 => x"08810580",
   123 => x"d6d40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480d6",
   128 => x"d8088105",
   129 => x"80d6d80c",
   130 => x"80d6d808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80d6d8",
   134 => x"0c80d6d4",
   135 => x"08810580",
   136 => x"d6d40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"d6dc0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"d6dc0c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280d6",
   177 => x"dc088407",
   178 => x"80d6dc0c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80d3",
   183 => x"8c0c8171",
   184 => x"2bff05f6",
   185 => x"880cfecc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80d6dc",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80d6",
   208 => x"c40c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"02dc050d",
  1093 => x"8059810b",
  1094 => x"ec0c840b",
  1095 => x"ec0c7a52",
  1096 => x"80d6e051",
  1097 => x"80c6fc2d",
  1098 => x"80d6c408",
  1099 => x"792e80f4",
  1100 => x"3880d6e4",
  1101 => x"0879ff12",
  1102 => x"56595673",
  1103 => x"792e8b38",
  1104 => x"81187481",
  1105 => x"2a555873",
  1106 => x"f738f718",
  1107 => x"58815980",
  1108 => x"762580d0",
  1109 => x"38775273",
  1110 => x"5184a82d",
  1111 => x"80d7b452",
  1112 => x"80d6e051",
  1113 => x"80c9d02d",
  1114 => x"80d6c408",
  1115 => x"802e9b38",
  1116 => x"80d7b457",
  1117 => x"83fc5576",
  1118 => x"70840558",
  1119 => x"08e80cfc",
  1120 => x"15557480",
  1121 => x"25f138a3",
  1122 => x"920480d6",
  1123 => x"c4085984",
  1124 => x"805680d6",
  1125 => x"e05180c9",
  1126 => x"9f2dfc80",
  1127 => x"16811555",
  1128 => x"56a2cf04",
  1129 => x"80d6e408",
  1130 => x"f80c8051",
  1131 => x"86da2d78",
  1132 => x"802e8838",
  1133 => x"80d39051",
  1134 => x"a3bf0480",
  1135 => x"d49451ab",
  1136 => x"b32d7880",
  1137 => x"d6c40c02",
  1138 => x"a4050d04",
  1139 => x"02f0050d",
  1140 => x"840bec0c",
  1141 => x"a8f02da5",
  1142 => x"a52d81f9",
  1143 => x"2d8352a8",
  1144 => x"d32d8151",
  1145 => x"858d2dff",
  1146 => x"12527180",
  1147 => x"25f13884",
  1148 => x"0bec0c80",
  1149 => x"d1c05186",
  1150 => x"a02dbdab",
  1151 => x"2d80d6c4",
  1152 => x"08802e81",
  1153 => x"8938a290",
  1154 => x"5180d0a5",
  1155 => x"2d80d390",
  1156 => x"51abb32d",
  1157 => x"a9922da5",
  1158 => x"b12dabc6",
  1159 => x"2d80d3a4",
  1160 => x"0b80f52d",
  1161 => x"80d58008",
  1162 => x"70810654",
  1163 => x"55537180",
  1164 => x"2e853872",
  1165 => x"84075373",
  1166 => x"812a7081",
  1167 => x"06515271",
  1168 => x"802e8538",
  1169 => x"72820753",
  1170 => x"73822a70",
  1171 => x"81065152",
  1172 => x"71802e85",
  1173 => x"38728107",
  1174 => x"5373832a",
  1175 => x"70810651",
  1176 => x"5271802e",
  1177 => x"85387288",
  1178 => x"07537384",
  1179 => x"2a708106",
  1180 => x"51527180",
  1181 => x"2e853872",
  1182 => x"90075372",
  1183 => x"fc0c8652",
  1184 => x"80d6c408",
  1185 => x"83388452",
  1186 => x"71ec0ca4",
  1187 => x"9704800b",
  1188 => x"80d6c40c",
  1189 => x"0290050d",
  1190 => x"0471980c",
  1191 => x"04ffb008",
  1192 => x"80d6c40c",
  1193 => x"04810bff",
  1194 => x"b00c0480",
  1195 => x"0bffb00c",
  1196 => x"0402f405",
  1197 => x"0da6bf04",
  1198 => x"80d6c408",
  1199 => x"81f02e09",
  1200 => x"81068a38",
  1201 => x"810b80d4",
  1202 => x"f80ca6bf",
  1203 => x"0480d6c4",
  1204 => x"0881e02e",
  1205 => x"0981068a",
  1206 => x"38810b80",
  1207 => x"d4fc0ca6",
  1208 => x"bf0480d6",
  1209 => x"c4085280",
  1210 => x"d4fc0880",
  1211 => x"2e893880",
  1212 => x"d6c40881",
  1213 => x"80055271",
  1214 => x"842c728f",
  1215 => x"06535380",
  1216 => x"d4f80880",
  1217 => x"2e9a3872",
  1218 => x"842980d4",
  1219 => x"b8057213",
  1220 => x"81712b70",
  1221 => x"09730806",
  1222 => x"730c5153",
  1223 => x"53a6b304",
  1224 => x"72842980",
  1225 => x"d4b80572",
  1226 => x"1383712b",
  1227 => x"72080772",
  1228 => x"0c535380",
  1229 => x"0b80d4fc",
  1230 => x"0c800b80",
  1231 => x"d4f80c80",
  1232 => x"d6ec51a7",
  1233 => x"c62d80d6",
  1234 => x"c408ff24",
  1235 => x"feea3880",
  1236 => x"0b80d6c4",
  1237 => x"0c028c05",
  1238 => x"0d0402f8",
  1239 => x"050d80d4",
  1240 => x"b8528f51",
  1241 => x"80727084",
  1242 => x"05540cff",
  1243 => x"11517080",
  1244 => x"25f23802",
  1245 => x"88050d04",
  1246 => x"02f0050d",
  1247 => x"7551a5ab",
  1248 => x"2d70822c",
  1249 => x"fc0680d4",
  1250 => x"b8117210",
  1251 => x"9e067108",
  1252 => x"70722a70",
  1253 => x"83068274",
  1254 => x"2b700974",
  1255 => x"06760c54",
  1256 => x"51565753",
  1257 => x"5153a5a5",
  1258 => x"2d7180d6",
  1259 => x"c40c0290",
  1260 => x"050d0402",
  1261 => x"fc050d72",
  1262 => x"5180710c",
  1263 => x"800b8412",
  1264 => x"0c028405",
  1265 => x"0d0402f0",
  1266 => x"050d7570",
  1267 => x"08841208",
  1268 => x"535353ff",
  1269 => x"5471712e",
  1270 => x"a838a5ab",
  1271 => x"2d841308",
  1272 => x"70842914",
  1273 => x"88117008",
  1274 => x"7081ff06",
  1275 => x"84180881",
  1276 => x"11870684",
  1277 => x"1a0c5351",
  1278 => x"55515151",
  1279 => x"a5a52d71",
  1280 => x"547380d6",
  1281 => x"c40c0290",
  1282 => x"050d0402",
  1283 => x"f8050da5",
  1284 => x"ab2de008",
  1285 => x"708b2a70",
  1286 => x"81065152",
  1287 => x"5270802e",
  1288 => x"a13880d6",
  1289 => x"ec087084",
  1290 => x"2980d6f4",
  1291 => x"057381ff",
  1292 => x"06710c51",
  1293 => x"5180d6ec",
  1294 => x"08811187",
  1295 => x"0680d6ec",
  1296 => x"0c51800b",
  1297 => x"80d7940c",
  1298 => x"a59d2da5",
  1299 => x"a52d0288",
  1300 => x"050d0402",
  1301 => x"fc050da5",
  1302 => x"ab2d810b",
  1303 => x"80d7940c",
  1304 => x"a5a52d80",
  1305 => x"d7940851",
  1306 => x"70f93802",
  1307 => x"84050d04",
  1308 => x"02fc050d",
  1309 => x"80d6ec51",
  1310 => x"a7b32da6",
  1311 => x"da2da88b",
  1312 => x"51a5992d",
  1313 => x"0284050d",
  1314 => x"0480d7a0",
  1315 => x"0880d6c4",
  1316 => x"0c0402fc",
  1317 => x"050d810b",
  1318 => x"80d5840c",
  1319 => x"8151858d",
  1320 => x"2d028405",
  1321 => x"0d0402fc",
  1322 => x"050da9b0",
  1323 => x"04a5b12d",
  1324 => x"80f651a6",
  1325 => x"f82d80d6",
  1326 => x"c408f238",
  1327 => x"80da51a6",
  1328 => x"f82d80d6",
  1329 => x"c408e638",
  1330 => x"80d6c408",
  1331 => x"80d5840c",
  1332 => x"80d6c408",
  1333 => x"51858d2d",
  1334 => x"0284050d",
  1335 => x"0402ec05",
  1336 => x"0d765480",
  1337 => x"52870b88",
  1338 => x"1580f52d",
  1339 => x"56537472",
  1340 => x"248338a0",
  1341 => x"53725183",
  1342 => x"842d8112",
  1343 => x"8b1580f5",
  1344 => x"2d545272",
  1345 => x"7225de38",
  1346 => x"0294050d",
  1347 => x"0402f005",
  1348 => x"0d80d7a0",
  1349 => x"085481f9",
  1350 => x"2d800b80",
  1351 => x"d7a40c73",
  1352 => x"08802e81",
  1353 => x"8938820b",
  1354 => x"80d6d80c",
  1355 => x"80d7a408",
  1356 => x"8f0680d6",
  1357 => x"d40c7308",
  1358 => x"5271832e",
  1359 => x"96387183",
  1360 => x"26893871",
  1361 => x"812eb038",
  1362 => x"ab970471",
  1363 => x"852ea038",
  1364 => x"ab970488",
  1365 => x"1480f52d",
  1366 => x"84150880",
  1367 => x"d1d85354",
  1368 => x"5286a02d",
  1369 => x"71842913",
  1370 => x"70085252",
  1371 => x"ab9b0473",
  1372 => x"51a9dd2d",
  1373 => x"ab970480",
  1374 => x"d5800888",
  1375 => x"15082c70",
  1376 => x"81065152",
  1377 => x"71802e88",
  1378 => x"3880d1dc",
  1379 => x"51ab9404",
  1380 => x"80d1e051",
  1381 => x"86a02d84",
  1382 => x"14085186",
  1383 => x"a02d80d7",
  1384 => x"a4088105",
  1385 => x"80d7a40c",
  1386 => x"8c1454aa",
  1387 => x"9f040290",
  1388 => x"050d0471",
  1389 => x"80d7a00c",
  1390 => x"aa8d2d80",
  1391 => x"d7a408ff",
  1392 => x"0580d7a8",
  1393 => x"0c0402e8",
  1394 => x"050d80d7",
  1395 => x"a00880d7",
  1396 => x"ac085755",
  1397 => x"80f651a6",
  1398 => x"f82d80d6",
  1399 => x"c408812a",
  1400 => x"70810651",
  1401 => x"5271802e",
  1402 => x"a438abf0",
  1403 => x"04a5b12d",
  1404 => x"80f651a6",
  1405 => x"f82d80d6",
  1406 => x"c408f238",
  1407 => x"80d58408",
  1408 => x"81327080",
  1409 => x"d5840c70",
  1410 => x"5252858d",
  1411 => x"2d800b80",
  1412 => x"d7980c80",
  1413 => x"0b80d79c",
  1414 => x"0c80d584",
  1415 => x"08838d38",
  1416 => x"80da51a6",
  1417 => x"f82d80d6",
  1418 => x"c408802e",
  1419 => x"8c3880d7",
  1420 => x"98088180",
  1421 => x"0780d798",
  1422 => x"0c80d951",
  1423 => x"a6f82d80",
  1424 => x"d6c40880",
  1425 => x"2e8c3880",
  1426 => x"d7980880",
  1427 => x"c00780d7",
  1428 => x"980c8194",
  1429 => x"51a6f82d",
  1430 => x"80d6c408",
  1431 => x"802e8b38",
  1432 => x"80d79808",
  1433 => x"900780d7",
  1434 => x"980c8191",
  1435 => x"51a6f82d",
  1436 => x"80d6c408",
  1437 => x"802e8b38",
  1438 => x"80d79808",
  1439 => x"a00780d7",
  1440 => x"980c81f5",
  1441 => x"51a6f82d",
  1442 => x"80d6c408",
  1443 => x"802e8b38",
  1444 => x"80d79808",
  1445 => x"810780d7",
  1446 => x"980c81f2",
  1447 => x"51a6f82d",
  1448 => x"80d6c408",
  1449 => x"802e8b38",
  1450 => x"80d79808",
  1451 => x"820780d7",
  1452 => x"980c81eb",
  1453 => x"51a6f82d",
  1454 => x"80d6c408",
  1455 => x"802e8b38",
  1456 => x"80d79808",
  1457 => x"840780d7",
  1458 => x"980c81f4",
  1459 => x"51a6f82d",
  1460 => x"80d6c408",
  1461 => x"802e8b38",
  1462 => x"80d79808",
  1463 => x"880780d7",
  1464 => x"980c80d8",
  1465 => x"51a6f82d",
  1466 => x"80d6c408",
  1467 => x"802e8c38",
  1468 => x"80d79c08",
  1469 => x"81800780",
  1470 => x"d79c0c92",
  1471 => x"51a6f82d",
  1472 => x"80d6c408",
  1473 => x"802e8c38",
  1474 => x"80d79c08",
  1475 => x"80c00780",
  1476 => x"d79c0c94",
  1477 => x"51a6f82d",
  1478 => x"80d6c408",
  1479 => x"802e8b38",
  1480 => x"80d79c08",
  1481 => x"900780d7",
  1482 => x"9c0c9151",
  1483 => x"a6f82d80",
  1484 => x"d6c40880",
  1485 => x"2e8b3880",
  1486 => x"d79c08a0",
  1487 => x"0780d79c",
  1488 => x"0c9d51a6",
  1489 => x"f82d80d6",
  1490 => x"c408802e",
  1491 => x"8b3880d7",
  1492 => x"9c088107",
  1493 => x"80d79c0c",
  1494 => x"9b51a6f8",
  1495 => x"2d80d6c4",
  1496 => x"08802e8b",
  1497 => x"3880d79c",
  1498 => x"08820780",
  1499 => x"d79c0c9c",
  1500 => x"51a6f82d",
  1501 => x"80d6c408",
  1502 => x"802e8b38",
  1503 => x"80d79c08",
  1504 => x"840780d7",
  1505 => x"9c0ca351",
  1506 => x"a6f82d80",
  1507 => x"d6c40880",
  1508 => x"2e8b3880",
  1509 => x"d79c0888",
  1510 => x"0780d79c",
  1511 => x"0c81fd51",
  1512 => x"a6f82d81",
  1513 => x"fa51a6f8",
  1514 => x"2db58104",
  1515 => x"81f551a6",
  1516 => x"f82d80d6",
  1517 => x"c408812a",
  1518 => x"70810651",
  1519 => x"5271802e",
  1520 => x"b33880d7",
  1521 => x"a8085271",
  1522 => x"802e8a38",
  1523 => x"ff1280d7",
  1524 => x"a80caff4",
  1525 => x"0480d7a4",
  1526 => x"081080d7",
  1527 => x"a4080570",
  1528 => x"84291651",
  1529 => x"52881208",
  1530 => x"802e8938",
  1531 => x"ff518812",
  1532 => x"0852712d",
  1533 => x"81f251a6",
  1534 => x"f82d80d6",
  1535 => x"c408812a",
  1536 => x"70810651",
  1537 => x"5271802e",
  1538 => x"b43880d7",
  1539 => x"a408ff11",
  1540 => x"80d7a808",
  1541 => x"56535373",
  1542 => x"72258a38",
  1543 => x"811480d7",
  1544 => x"a80cb0bd",
  1545 => x"04721013",
  1546 => x"70842916",
  1547 => x"51528812",
  1548 => x"08802e89",
  1549 => x"38fe5188",
  1550 => x"12085271",
  1551 => x"2d81fd51",
  1552 => x"a6f82d80",
  1553 => x"d6c40881",
  1554 => x"2a708106",
  1555 => x"51527180",
  1556 => x"2eb13880",
  1557 => x"d7a80880",
  1558 => x"2e8a3880",
  1559 => x"0b80d7a8",
  1560 => x"0cb18304",
  1561 => x"80d7a408",
  1562 => x"1080d7a4",
  1563 => x"08057084",
  1564 => x"29165152",
  1565 => x"88120880",
  1566 => x"2e8938fd",
  1567 => x"51881208",
  1568 => x"52712d81",
  1569 => x"fa51a6f8",
  1570 => x"2d80d6c4",
  1571 => x"08812a70",
  1572 => x"81065152",
  1573 => x"71802eb1",
  1574 => x"3880d7a4",
  1575 => x"08ff1154",
  1576 => x"5280d7a8",
  1577 => x"08732589",
  1578 => x"387280d7",
  1579 => x"a80cb1c9",
  1580 => x"04711012",
  1581 => x"70842916",
  1582 => x"51528812",
  1583 => x"08802e89",
  1584 => x"38fc5188",
  1585 => x"12085271",
  1586 => x"2d80d7a8",
  1587 => x"08705354",
  1588 => x"73802e8a",
  1589 => x"388c15ff",
  1590 => x"155555b1",
  1591 => x"d004820b",
  1592 => x"80d6d80c",
  1593 => x"718f0680",
  1594 => x"d6d40c81",
  1595 => x"eb51a6f8",
  1596 => x"2d80d6c4",
  1597 => x"08812a70",
  1598 => x"81065152",
  1599 => x"71802ead",
  1600 => x"38740885",
  1601 => x"2e098106",
  1602 => x"a4388815",
  1603 => x"80f52dff",
  1604 => x"05527188",
  1605 => x"1681b72d",
  1606 => x"71982b52",
  1607 => x"71802588",
  1608 => x"38800b88",
  1609 => x"1681b72d",
  1610 => x"7451a9dd",
  1611 => x"2d81f451",
  1612 => x"a6f82d80",
  1613 => x"d6c40881",
  1614 => x"2a708106",
  1615 => x"51527180",
  1616 => x"2eb33874",
  1617 => x"08852e09",
  1618 => x"8106aa38",
  1619 => x"881580f5",
  1620 => x"2d810552",
  1621 => x"71881681",
  1622 => x"b72d7181",
  1623 => x"ff068b16",
  1624 => x"80f52d54",
  1625 => x"52727227",
  1626 => x"87387288",
  1627 => x"1681b72d",
  1628 => x"7451a9dd",
  1629 => x"2d80da51",
  1630 => x"a6f82d80",
  1631 => x"d6c40881",
  1632 => x"2a708106",
  1633 => x"51527180",
  1634 => x"2e81ad38",
  1635 => x"80d7a008",
  1636 => x"80d7a808",
  1637 => x"55537380",
  1638 => x"2e8a388c",
  1639 => x"13ff1555",
  1640 => x"53b39604",
  1641 => x"72085271",
  1642 => x"822ea638",
  1643 => x"71822689",
  1644 => x"3871812e",
  1645 => x"aa38b4b8",
  1646 => x"0471832e",
  1647 => x"b4387184",
  1648 => x"2e098106",
  1649 => x"80f23888",
  1650 => x"130851ab",
  1651 => x"b32db4b8",
  1652 => x"0480d7a8",
  1653 => x"08518813",
  1654 => x"0852712d",
  1655 => x"b4b80481",
  1656 => x"0b881408",
  1657 => x"2b80d580",
  1658 => x"083280d5",
  1659 => x"800cb48c",
  1660 => x"04881380",
  1661 => x"f52d8105",
  1662 => x"8b1480f5",
  1663 => x"2d535471",
  1664 => x"74248338",
  1665 => x"80547388",
  1666 => x"1481b72d",
  1667 => x"aa8d2db4",
  1668 => x"b8047508",
  1669 => x"802ea438",
  1670 => x"750851a6",
  1671 => x"f82d80d6",
  1672 => x"c4088106",
  1673 => x"5271802e",
  1674 => x"8c3880d7",
  1675 => x"a8085184",
  1676 => x"16085271",
  1677 => x"2d881656",
  1678 => x"75d83880",
  1679 => x"54800b80",
  1680 => x"d6d80c73",
  1681 => x"8f0680d6",
  1682 => x"d40ca052",
  1683 => x"7380d7a8",
  1684 => x"082e0981",
  1685 => x"06993880",
  1686 => x"d7a408ff",
  1687 => x"05743270",
  1688 => x"09810570",
  1689 => x"72079f2a",
  1690 => x"91713151",
  1691 => x"51535371",
  1692 => x"5183842d",
  1693 => x"8114548e",
  1694 => x"7425c238",
  1695 => x"80d58408",
  1696 => x"527180d6",
  1697 => x"c40c0298",
  1698 => x"050d0402",
  1699 => x"f4050dd4",
  1700 => x"5281ff72",
  1701 => x"0c710853",
  1702 => x"81ff720c",
  1703 => x"72882b83",
  1704 => x"fe800672",
  1705 => x"087081ff",
  1706 => x"06515253",
  1707 => x"81ff720c",
  1708 => x"72710788",
  1709 => x"2b720870",
  1710 => x"81ff0651",
  1711 => x"525381ff",
  1712 => x"720c7271",
  1713 => x"07882b72",
  1714 => x"087081ff",
  1715 => x"06720780",
  1716 => x"d6c40c52",
  1717 => x"53028c05",
  1718 => x"0d0402f4",
  1719 => x"050d7476",
  1720 => x"7181ff06",
  1721 => x"d40c5353",
  1722 => x"80d7b008",
  1723 => x"85387189",
  1724 => x"2b527198",
  1725 => x"2ad40c71",
  1726 => x"902a7081",
  1727 => x"ff06d40c",
  1728 => x"5171882a",
  1729 => x"7081ff06",
  1730 => x"d40c5171",
  1731 => x"81ff06d4",
  1732 => x"0c72902a",
  1733 => x"7081ff06",
  1734 => x"d40c51d4",
  1735 => x"087081ff",
  1736 => x"06515182",
  1737 => x"b8bf5270",
  1738 => x"81ff2e09",
  1739 => x"81069438",
  1740 => x"81ff0bd4",
  1741 => x"0cd40870",
  1742 => x"81ff06ff",
  1743 => x"14545151",
  1744 => x"71e53870",
  1745 => x"80d6c40c",
  1746 => x"028c050d",
  1747 => x"0402fc05",
  1748 => x"0d81c751",
  1749 => x"81ff0bd4",
  1750 => x"0cff1151",
  1751 => x"708025f4",
  1752 => x"38028405",
  1753 => x"0d0402f4",
  1754 => x"050d81ff",
  1755 => x"0bd40c93",
  1756 => x"53805287",
  1757 => x"fc80c151",
  1758 => x"b5da2d80",
  1759 => x"d6c4088b",
  1760 => x"3881ff0b",
  1761 => x"d40c8153",
  1762 => x"b79404b6",
  1763 => x"cd2dff13",
  1764 => x"5372de38",
  1765 => x"7280d6c4",
  1766 => x"0c028c05",
  1767 => x"0d0402ec",
  1768 => x"050d810b",
  1769 => x"80d7b00c",
  1770 => x"8454d008",
  1771 => x"708f2a70",
  1772 => x"81065151",
  1773 => x"5372f338",
  1774 => x"72d00cb6",
  1775 => x"cd2d80d1",
  1776 => x"e45186a0",
  1777 => x"2dd00870",
  1778 => x"8f2a7081",
  1779 => x"06515153",
  1780 => x"72f33881",
  1781 => x"0bd00cb1",
  1782 => x"53805284",
  1783 => x"d480c051",
  1784 => x"b5da2d80",
  1785 => x"d6c40881",
  1786 => x"2e933872",
  1787 => x"822ebf38",
  1788 => x"ff135372",
  1789 => x"e438ff14",
  1790 => x"5473ffae",
  1791 => x"38b6cd2d",
  1792 => x"83aa5284",
  1793 => x"9c80c851",
  1794 => x"b5da2d80",
  1795 => x"d6c40881",
  1796 => x"2e098106",
  1797 => x"9338b58b",
  1798 => x"2d80d6c4",
  1799 => x"0883ffff",
  1800 => x"06537283",
  1801 => x"aa2e9f38",
  1802 => x"b6e62db8",
  1803 => x"c10480d1",
  1804 => x"f05186a0",
  1805 => x"2d8053ba",
  1806 => x"960480d2",
  1807 => x"885186a0",
  1808 => x"2d8054b9",
  1809 => x"e70481ff",
  1810 => x"0bd40cb1",
  1811 => x"54b6cd2d",
  1812 => x"8fcf5380",
  1813 => x"5287fc80",
  1814 => x"f751b5da",
  1815 => x"2d80d6c4",
  1816 => x"085580d6",
  1817 => x"c408812e",
  1818 => x"0981069c",
  1819 => x"3881ff0b",
  1820 => x"d40c820a",
  1821 => x"52849c80",
  1822 => x"e951b5da",
  1823 => x"2d80d6c4",
  1824 => x"08802e8d",
  1825 => x"38b6cd2d",
  1826 => x"ff135372",
  1827 => x"c638b9da",
  1828 => x"0481ff0b",
  1829 => x"d40c80d6",
  1830 => x"c4085287",
  1831 => x"fc80fa51",
  1832 => x"b5da2d80",
  1833 => x"d6c408b2",
  1834 => x"3881ff0b",
  1835 => x"d40cd408",
  1836 => x"5381ff0b",
  1837 => x"d40c81ff",
  1838 => x"0bd40c81",
  1839 => x"ff0bd40c",
  1840 => x"81ff0bd4",
  1841 => x"0c72862a",
  1842 => x"70810676",
  1843 => x"56515372",
  1844 => x"963880d6",
  1845 => x"c40854b9",
  1846 => x"e7047382",
  1847 => x"2efedb38",
  1848 => x"ff145473",
  1849 => x"fee73873",
  1850 => x"80d7b00c",
  1851 => x"738b3881",
  1852 => x"5287fc80",
  1853 => x"d051b5da",
  1854 => x"2d81ff0b",
  1855 => x"d40cd008",
  1856 => x"708f2a70",
  1857 => x"81065151",
  1858 => x"5372f338",
  1859 => x"72d00c81",
  1860 => x"ff0bd40c",
  1861 => x"81537280",
  1862 => x"d6c40c02",
  1863 => x"94050d04",
  1864 => x"02e8050d",
  1865 => x"78558056",
  1866 => x"81ff0bd4",
  1867 => x"0cd00870",
  1868 => x"8f2a7081",
  1869 => x"06515153",
  1870 => x"72f33882",
  1871 => x"810bd00c",
  1872 => x"81ff0bd4",
  1873 => x"0c775287",
  1874 => x"fc80d151",
  1875 => x"b5da2d80",
  1876 => x"dbc6df54",
  1877 => x"80d6c408",
  1878 => x"802e8b38",
  1879 => x"80d2a851",
  1880 => x"86a02dbb",
  1881 => x"ba0481ff",
  1882 => x"0bd40cd4",
  1883 => x"087081ff",
  1884 => x"06515372",
  1885 => x"81fe2e09",
  1886 => x"81069e38",
  1887 => x"80ff53b5",
  1888 => x"8b2d80d6",
  1889 => x"c4087570",
  1890 => x"8405570c",
  1891 => x"ff135372",
  1892 => x"8025ec38",
  1893 => x"8156bb9f",
  1894 => x"04ff1454",
  1895 => x"73c83881",
  1896 => x"ff0bd40c",
  1897 => x"81ff0bd4",
  1898 => x"0cd00870",
  1899 => x"8f2a7081",
  1900 => x"06515153",
  1901 => x"72f33872",
  1902 => x"d00c7580",
  1903 => x"d6c40c02",
  1904 => x"98050d04",
  1905 => x"02e8050d",
  1906 => x"77797b58",
  1907 => x"55558053",
  1908 => x"727625a3",
  1909 => x"38747081",
  1910 => x"055680f5",
  1911 => x"2d747081",
  1912 => x"055680f5",
  1913 => x"2d525271",
  1914 => x"712e8638",
  1915 => x"8151bbf9",
  1916 => x"04811353",
  1917 => x"bbd00480",
  1918 => x"517080d6",
  1919 => x"c40c0298",
  1920 => x"050d0402",
  1921 => x"ec050d76",
  1922 => x"5574802e",
  1923 => x"80c4389a",
  1924 => x"1580e02d",
  1925 => x"5180caaa",
  1926 => x"2d80d6c4",
  1927 => x"0880d6c4",
  1928 => x"0880dde4",
  1929 => x"0c80d6c4",
  1930 => x"08545480",
  1931 => x"ddc00880",
  1932 => x"2e9b3894",
  1933 => x"1580e02d",
  1934 => x"5180caaa",
  1935 => x"2d80d6c4",
  1936 => x"08902b83",
  1937 => x"fff00a06",
  1938 => x"70750751",
  1939 => x"537280dd",
  1940 => x"e40c80dd",
  1941 => x"e4085372",
  1942 => x"802e9d38",
  1943 => x"80ddb808",
  1944 => x"fe147129",
  1945 => x"80ddcc08",
  1946 => x"0580dde8",
  1947 => x"0c70842b",
  1948 => x"80ddc40c",
  1949 => x"54bda604",
  1950 => x"80ddd008",
  1951 => x"80dde40c",
  1952 => x"80ddd408",
  1953 => x"80dde80c",
  1954 => x"80ddc008",
  1955 => x"802e8b38",
  1956 => x"80ddb808",
  1957 => x"842b53bd",
  1958 => x"a10480dd",
  1959 => x"d808842b",
  1960 => x"537280dd",
  1961 => x"c40c0294",
  1962 => x"050d0402",
  1963 => x"d8050d80",
  1964 => x"0b80ddc0",
  1965 => x"0c8454b7",
  1966 => x"9e2d80d6",
  1967 => x"c408802e",
  1968 => x"973880d7",
  1969 => x"b4528051",
  1970 => x"baa02d80",
  1971 => x"d6c40880",
  1972 => x"2e8638fe",
  1973 => x"54bde004",
  1974 => x"ff145473",
  1975 => x"8024d838",
  1976 => x"738e3880",
  1977 => x"d2b85186",
  1978 => x"a02d7355",
  1979 => x"80c3ba04",
  1980 => x"8056810b",
  1981 => x"80ddec0c",
  1982 => x"885380d2",
  1983 => x"cc5280d7",
  1984 => x"ea51bbc4",
  1985 => x"2d80d6c4",
  1986 => x"08762e09",
  1987 => x"81068938",
  1988 => x"80d6c408",
  1989 => x"80ddec0c",
  1990 => x"885380d2",
  1991 => x"d85280d8",
  1992 => x"8651bbc4",
  1993 => x"2d80d6c4",
  1994 => x"08893880",
  1995 => x"d6c40880",
  1996 => x"ddec0c80",
  1997 => x"ddec0880",
  1998 => x"2e818238",
  1999 => x"80dafa0b",
  2000 => x"80f52d80",
  2001 => x"dafb0b80",
  2002 => x"f52d7198",
  2003 => x"2b71902b",
  2004 => x"0780dafc",
  2005 => x"0b80f52d",
  2006 => x"70882b72",
  2007 => x"0780dafd",
  2008 => x"0b80f52d",
  2009 => x"710780db",
  2010 => x"b20b80f5",
  2011 => x"2d80dbb3",
  2012 => x"0b80f52d",
  2013 => x"71882b07",
  2014 => x"535f5452",
  2015 => x"5a565755",
  2016 => x"7381abaa",
  2017 => x"2e098106",
  2018 => x"8f387551",
  2019 => x"80c9f92d",
  2020 => x"80d6c408",
  2021 => x"56bfa604",
  2022 => x"7382d4d5",
  2023 => x"2e883880",
  2024 => x"d2e451bf",
  2025 => x"f20480d7",
  2026 => x"b4527551",
  2027 => x"baa02d80",
  2028 => x"d6c40855",
  2029 => x"80d6c408",
  2030 => x"802e83fe",
  2031 => x"38885380",
  2032 => x"d2d85280",
  2033 => x"d88651bb",
  2034 => x"c42d80d6",
  2035 => x"c4088a38",
  2036 => x"810b80dd",
  2037 => x"c00cbff9",
  2038 => x"04885380",
  2039 => x"d2cc5280",
  2040 => x"d7ea51bb",
  2041 => x"c42d80d6",
  2042 => x"c408802e",
  2043 => x"8c3880d2",
  2044 => x"f85186a0",
  2045 => x"2d80c0d8",
  2046 => x"0480dbb2",
  2047 => x"0b80f52d",
  2048 => x"547380d5",
  2049 => x"2e098106",
  2050 => x"80ce3880",
  2051 => x"dbb30b80",
  2052 => x"f52d5473",
  2053 => x"81aa2e09",
  2054 => x"8106bd38",
  2055 => x"800b80d7",
  2056 => x"b40b80f5",
  2057 => x"2d565474",
  2058 => x"81e92e83",
  2059 => x"38815474",
  2060 => x"81eb2e8c",
  2061 => x"38805573",
  2062 => x"752e0981",
  2063 => x"0682fb38",
  2064 => x"80d7bf0b",
  2065 => x"80f52d55",
  2066 => x"748e3880",
  2067 => x"d7c00b80",
  2068 => x"f52d5473",
  2069 => x"822e8738",
  2070 => x"805580c3",
  2071 => x"ba0480d7",
  2072 => x"c10b80f5",
  2073 => x"2d7080dd",
  2074 => x"b80cff05",
  2075 => x"80ddbc0c",
  2076 => x"80d7c20b",
  2077 => x"80f52d80",
  2078 => x"d7c30b80",
  2079 => x"f52d5876",
  2080 => x"05778280",
  2081 => x"29057080",
  2082 => x"ddc80c80",
  2083 => x"d7c40b80",
  2084 => x"f52d7080",
  2085 => x"dddc0c80",
  2086 => x"ddc00859",
  2087 => x"57587680",
  2088 => x"2e81b838",
  2089 => x"885380d2",
  2090 => x"d85280d8",
  2091 => x"8651bbc4",
  2092 => x"2d80d6c4",
  2093 => x"08828338",
  2094 => x"80ddb808",
  2095 => x"70842b80",
  2096 => x"ddc40c70",
  2097 => x"80ddd80c",
  2098 => x"80d7d90b",
  2099 => x"80f52d80",
  2100 => x"d7d80b80",
  2101 => x"f52d7182",
  2102 => x"80290580",
  2103 => x"d7da0b80",
  2104 => x"f52d7084",
  2105 => x"80802912",
  2106 => x"80d7db0b",
  2107 => x"80f52d70",
  2108 => x"81800a29",
  2109 => x"127080dd",
  2110 => x"e00c80dd",
  2111 => x"dc087129",
  2112 => x"80ddc808",
  2113 => x"057080dd",
  2114 => x"cc0c80d7",
  2115 => x"e10b80f5",
  2116 => x"2d80d7e0",
  2117 => x"0b80f52d",
  2118 => x"71828029",
  2119 => x"0580d7e2",
  2120 => x"0b80f52d",
  2121 => x"70848080",
  2122 => x"291280d7",
  2123 => x"e30b80f5",
  2124 => x"2d70982b",
  2125 => x"81f00a06",
  2126 => x"72057080",
  2127 => x"ddd00cfe",
  2128 => x"117e2977",
  2129 => x"0580ddd4",
  2130 => x"0c525952",
  2131 => x"43545e51",
  2132 => x"5259525d",
  2133 => x"57595780",
  2134 => x"c3b30480",
  2135 => x"d7c60b80",
  2136 => x"f52d80d7",
  2137 => x"c50b80f5",
  2138 => x"2d718280",
  2139 => x"29057080",
  2140 => x"ddc40c70",
  2141 => x"a02983ff",
  2142 => x"0570892a",
  2143 => x"7080ddd8",
  2144 => x"0c80d7cb",
  2145 => x"0b80f52d",
  2146 => x"80d7ca0b",
  2147 => x"80f52d71",
  2148 => x"82802905",
  2149 => x"7080dde0",
  2150 => x"0c7b7129",
  2151 => x"1e7080dd",
  2152 => x"d40c7d80",
  2153 => x"ddd00c73",
  2154 => x"0580ddcc",
  2155 => x"0c555e51",
  2156 => x"51555580",
  2157 => x"51bc832d",
  2158 => x"81557480",
  2159 => x"d6c40c02",
  2160 => x"a8050d04",
  2161 => x"02ec050d",
  2162 => x"7670872c",
  2163 => x"7180ff06",
  2164 => x"55565480",
  2165 => x"ddc0088a",
  2166 => x"3873882c",
  2167 => x"7481ff06",
  2168 => x"545580d7",
  2169 => x"b45280dd",
  2170 => x"c8081551",
  2171 => x"baa02d80",
  2172 => x"d6c40854",
  2173 => x"80d6c408",
  2174 => x"802ebb38",
  2175 => x"80ddc008",
  2176 => x"802e9c38",
  2177 => x"72842980",
  2178 => x"d7b40570",
  2179 => x"08525380",
  2180 => x"c9f92d80",
  2181 => x"d6c408f0",
  2182 => x"0a065380",
  2183 => x"c4b40472",
  2184 => x"1080d7b4",
  2185 => x"057080e0",
  2186 => x"2d525380",
  2187 => x"caaa2d80",
  2188 => x"d6c40853",
  2189 => x"72547380",
  2190 => x"d6c40c02",
  2191 => x"94050d04",
  2192 => x"02e0050d",
  2193 => x"7970842c",
  2194 => x"80dde808",
  2195 => x"05718f06",
  2196 => x"52555372",
  2197 => x"8a3880d7",
  2198 => x"b4527351",
  2199 => x"baa02d72",
  2200 => x"a02980d7",
  2201 => x"b4055480",
  2202 => x"7480f52d",
  2203 => x"56537473",
  2204 => x"2e833881",
  2205 => x"537481e5",
  2206 => x"2e81f538",
  2207 => x"81707406",
  2208 => x"54587280",
  2209 => x"2e81e938",
  2210 => x"8b1480f5",
  2211 => x"2d70832a",
  2212 => x"79065856",
  2213 => x"769c3880",
  2214 => x"d5880853",
  2215 => x"72893872",
  2216 => x"80dbb40b",
  2217 => x"81b72d76",
  2218 => x"80d5880c",
  2219 => x"735380c6",
  2220 => x"f204758f",
  2221 => x"2e098106",
  2222 => x"81b63874",
  2223 => x"9f068d29",
  2224 => x"80dba711",
  2225 => x"51538114",
  2226 => x"80f52d73",
  2227 => x"70810555",
  2228 => x"81b72d83",
  2229 => x"1480f52d",
  2230 => x"73708105",
  2231 => x"5581b72d",
  2232 => x"851480f5",
  2233 => x"2d737081",
  2234 => x"055581b7",
  2235 => x"2d871480",
  2236 => x"f52d7370",
  2237 => x"81055581",
  2238 => x"b72d8914",
  2239 => x"80f52d73",
  2240 => x"70810555",
  2241 => x"81b72d8e",
  2242 => x"1480f52d",
  2243 => x"73708105",
  2244 => x"5581b72d",
  2245 => x"901480f5",
  2246 => x"2d737081",
  2247 => x"055581b7",
  2248 => x"2d921480",
  2249 => x"f52d7370",
  2250 => x"81055581",
  2251 => x"b72d9414",
  2252 => x"80f52d73",
  2253 => x"70810555",
  2254 => x"81b72d96",
  2255 => x"1480f52d",
  2256 => x"73708105",
  2257 => x"5581b72d",
  2258 => x"981480f5",
  2259 => x"2d737081",
  2260 => x"055581b7",
  2261 => x"2d9c1480",
  2262 => x"f52d7370",
  2263 => x"81055581",
  2264 => x"b72d9e14",
  2265 => x"80f52d73",
  2266 => x"81b72d77",
  2267 => x"80d5880c",
  2268 => x"80537280",
  2269 => x"d6c40c02",
  2270 => x"a0050d04",
  2271 => x"02cc050d",
  2272 => x"7e605e5a",
  2273 => x"800b80dd",
  2274 => x"e40880dd",
  2275 => x"e808595c",
  2276 => x"56805880",
  2277 => x"ddc40878",
  2278 => x"2e81bc38",
  2279 => x"778f06a0",
  2280 => x"17575473",
  2281 => x"913880d7",
  2282 => x"b4527651",
  2283 => x"811757ba",
  2284 => x"a02d80d7",
  2285 => x"b4568076",
  2286 => x"80f52d56",
  2287 => x"5474742e",
  2288 => x"83388154",
  2289 => x"7481e52e",
  2290 => x"81813881",
  2291 => x"70750655",
  2292 => x"5c73802e",
  2293 => x"80f5388b",
  2294 => x"1680f52d",
  2295 => x"98065978",
  2296 => x"80e9388b",
  2297 => x"537c5275",
  2298 => x"51bbc42d",
  2299 => x"80d6c408",
  2300 => x"80d9389c",
  2301 => x"16085180",
  2302 => x"c9f92d80",
  2303 => x"d6c40884",
  2304 => x"1b0c9a16",
  2305 => x"80e02d51",
  2306 => x"80caaa2d",
  2307 => x"80d6c408",
  2308 => x"80d6c408",
  2309 => x"881c0c80",
  2310 => x"d6c40855",
  2311 => x"5580ddc0",
  2312 => x"08802e9a",
  2313 => x"38941680",
  2314 => x"e02d5180",
  2315 => x"caaa2d80",
  2316 => x"d6c40890",
  2317 => x"2b83fff0",
  2318 => x"0a067016",
  2319 => x"51547388",
  2320 => x"1b0c787a",
  2321 => x"0c7b5480",
  2322 => x"c9950481",
  2323 => x"185880dd",
  2324 => x"c4087826",
  2325 => x"fec63880",
  2326 => x"ddc00880",
  2327 => x"2eb5387a",
  2328 => x"5180c3c4",
  2329 => x"2d80d6c4",
  2330 => x"0880d6c4",
  2331 => x"0880ffff",
  2332 => x"fff80655",
  2333 => x"5b7380ff",
  2334 => x"fffff82e",
  2335 => x"963880d6",
  2336 => x"c408fe05",
  2337 => x"80ddb808",
  2338 => x"2980ddcc",
  2339 => x"08055780",
  2340 => x"c7910480",
  2341 => x"547380d6",
  2342 => x"c40c02b4",
  2343 => x"050d0402",
  2344 => x"f4050d74",
  2345 => x"70088105",
  2346 => x"710c7008",
  2347 => x"80ddbc08",
  2348 => x"06535371",
  2349 => x"90388813",
  2350 => x"085180c3",
  2351 => x"c42d80d6",
  2352 => x"c4088814",
  2353 => x"0c810b80",
  2354 => x"d6c40c02",
  2355 => x"8c050d04",
  2356 => x"02f0050d",
  2357 => x"75881108",
  2358 => x"fe0580dd",
  2359 => x"b8082980",
  2360 => x"ddcc0811",
  2361 => x"720880dd",
  2362 => x"bc080605",
  2363 => x"79555354",
  2364 => x"54baa02d",
  2365 => x"0290050d",
  2366 => x"0402f405",
  2367 => x"0d747088",
  2368 => x"2a83fe80",
  2369 => x"06707298",
  2370 => x"2a077288",
  2371 => x"2b87fc80",
  2372 => x"80067398",
  2373 => x"2b81f00a",
  2374 => x"06717307",
  2375 => x"0780d6c4",
  2376 => x"0c565153",
  2377 => x"51028c05",
  2378 => x"0d0402f8",
  2379 => x"050d028e",
  2380 => x"0580f52d",
  2381 => x"74882b07",
  2382 => x"7083ffff",
  2383 => x"0680d6c4",
  2384 => x"0c510288",
  2385 => x"050d0402",
  2386 => x"f4050d74",
  2387 => x"76785354",
  2388 => x"52807125",
  2389 => x"97387270",
  2390 => x"81055480",
  2391 => x"f52d7270",
  2392 => x"81055481",
  2393 => x"b72dff11",
  2394 => x"5170eb38",
  2395 => x"807281b7",
  2396 => x"2d028c05",
  2397 => x"0d0402e8",
  2398 => x"050d7756",
  2399 => x"80705654",
  2400 => x"737624b7",
  2401 => x"3880ddc4",
  2402 => x"08742eaf",
  2403 => x"38735180",
  2404 => x"c4c02d80",
  2405 => x"d6c40880",
  2406 => x"d6c40809",
  2407 => x"81057080",
  2408 => x"d6c40807",
  2409 => x"9f2a7705",
  2410 => x"81175757",
  2411 => x"53537476",
  2412 => x"24893880",
  2413 => x"ddc40874",
  2414 => x"26d33872",
  2415 => x"80d6c40c",
  2416 => x"0298050d",
  2417 => x"0402f005",
  2418 => x"0d80d6c0",
  2419 => x"08165180",
  2420 => x"caf62d80",
  2421 => x"d6c40880",
  2422 => x"2ea0388b",
  2423 => x"5380d6c4",
  2424 => x"085280db",
  2425 => x"b45180ca",
  2426 => x"c72d80dd",
  2427 => x"f0085473",
  2428 => x"802e8738",
  2429 => x"80dbb451",
  2430 => x"732d0290",
  2431 => x"050d0402",
  2432 => x"dc050d80",
  2433 => x"705a5574",
  2434 => x"80d6c008",
  2435 => x"25b53880",
  2436 => x"ddc40875",
  2437 => x"2ead3878",
  2438 => x"5180c4c0",
  2439 => x"2d80d6c4",
  2440 => x"08098105",
  2441 => x"7080d6c4",
  2442 => x"08079f2a",
  2443 => x"7605811b",
  2444 => x"5b565474",
  2445 => x"80d6c008",
  2446 => x"25893880",
  2447 => x"ddc40879",
  2448 => x"26d53880",
  2449 => x"557880dd",
  2450 => x"c4082781",
  2451 => x"e4387851",
  2452 => x"80c4c02d",
  2453 => x"80d6c408",
  2454 => x"802e81b4",
  2455 => x"3880d6c4",
  2456 => x"088b0580",
  2457 => x"f52d7084",
  2458 => x"2a708106",
  2459 => x"77107884",
  2460 => x"2b80dbb4",
  2461 => x"0b80f52d",
  2462 => x"5c5c5351",
  2463 => x"55567380",
  2464 => x"2e80ce38",
  2465 => x"7416822b",
  2466 => x"80ced50b",
  2467 => x"80d59412",
  2468 => x"0c547775",
  2469 => x"311080dd",
  2470 => x"f4115556",
  2471 => x"90747081",
  2472 => x"055681b7",
  2473 => x"2da07481",
  2474 => x"b72d7681",
  2475 => x"ff068116",
  2476 => x"58547380",
  2477 => x"2e8b389c",
  2478 => x"5380dbb4",
  2479 => x"5280cdc8",
  2480 => x"048b5380",
  2481 => x"d6c40852",
  2482 => x"80ddf616",
  2483 => x"5180ce86",
  2484 => x"04741682",
  2485 => x"2b80cbc5",
  2486 => x"0b80d594",
  2487 => x"120c5476",
  2488 => x"81ff0681",
  2489 => x"16585473",
  2490 => x"802e8b38",
  2491 => x"9c5380db",
  2492 => x"b45280cd",
  2493 => x"fd048b53",
  2494 => x"80d6c408",
  2495 => x"52777531",
  2496 => x"1080ddf4",
  2497 => x"05517655",
  2498 => x"80cac72d",
  2499 => x"80cea504",
  2500 => x"74902975",
  2501 => x"31701080",
  2502 => x"ddf40551",
  2503 => x"5480d6c4",
  2504 => x"087481b7",
  2505 => x"2d811959",
  2506 => x"748b24a4",
  2507 => x"3880ccc5",
  2508 => x"04749029",
  2509 => x"75317010",
  2510 => x"80ddf405",
  2511 => x"8c773157",
  2512 => x"51548074",
  2513 => x"81b72d9e",
  2514 => x"14ff1656",
  2515 => x"5474f338",
  2516 => x"02a4050d",
  2517 => x"0402fc05",
  2518 => x"0d80d6c0",
  2519 => x"08135180",
  2520 => x"caf62d80",
  2521 => x"d6c40880",
  2522 => x"2e893880",
  2523 => x"d6c40851",
  2524 => x"bc832d80",
  2525 => x"0b80d6c0",
  2526 => x"0c80cbff",
  2527 => x"2daa8d2d",
  2528 => x"0284050d",
  2529 => x"0402fc05",
  2530 => x"0d725170",
  2531 => x"fd2eb238",
  2532 => x"70fd248b",
  2533 => x"3870fc2e",
  2534 => x"80d03880",
  2535 => x"cff40470",
  2536 => x"fe2eb938",
  2537 => x"70ff2e09",
  2538 => x"810680c8",
  2539 => x"3880d6c0",
  2540 => x"08517080",
  2541 => x"2ebe38ff",
  2542 => x"1180d6c0",
  2543 => x"0c80cff4",
  2544 => x"0480d6c0",
  2545 => x"08f00570",
  2546 => x"80d6c00c",
  2547 => x"51708025",
  2548 => x"a338800b",
  2549 => x"80d6c00c",
  2550 => x"80cff404",
  2551 => x"80d6c008",
  2552 => x"810580d6",
  2553 => x"c00c80cf",
  2554 => x"f40480d6",
  2555 => x"c0089005",
  2556 => x"80d6c00c",
  2557 => x"80cbff2d",
  2558 => x"aa8d2d02",
  2559 => x"84050d04",
  2560 => x"02fc050d",
  2561 => x"800b80d6",
  2562 => x"c00c80cb",
  2563 => x"ff2da989",
  2564 => x"2d80d6c4",
  2565 => x"0880d6b0",
  2566 => x"0c80d58c",
  2567 => x"51abb32d",
  2568 => x"0284050d",
  2569 => x"047180dd",
  2570 => x"f00c0400",
  2571 => x"00ffffff",
  2572 => x"ff00ffff",
  2573 => x"ffff00ff",
  2574 => x"ffffff00",
  2575 => x"52657365",
  2576 => x"74000000",
  2577 => x"5363616e",
  2578 => x"6c696e65",
  2579 => x"73000000",
  2580 => x"50414c20",
  2581 => x"2f204e54",
  2582 => x"53430000",
  2583 => x"436f6c6f",
  2584 => x"72000000",
  2585 => x"44696666",
  2586 => x"6963756c",
  2587 => x"74792041",
  2588 => x"00000000",
  2589 => x"44696666",
  2590 => x"6963756c",
  2591 => x"74792042",
  2592 => x"00000000",
  2593 => x"53656c65",
  2594 => x"63740000",
  2595 => x"53746172",
  2596 => x"74000000",
  2597 => x"4c6f6164",
  2598 => x"20524f4d",
  2599 => x"20100000",
  2600 => x"45786974",
  2601 => x"00000000",
  2602 => x"524f4d20",
  2603 => x"6c6f6164",
  2604 => x"696e6720",
  2605 => x"6661696c",
  2606 => x"65640000",
  2607 => x"4f4b0000",
  2608 => x"496e6974",
  2609 => x"69616c69",
  2610 => x"7a696e67",
  2611 => x"20534420",
  2612 => x"63617264",
  2613 => x"0a000000",
  2614 => x"16200000",
  2615 => x"14200000",
  2616 => x"15200000",
  2617 => x"53442069",
  2618 => x"6e69742e",
  2619 => x"2e2e0a00",
  2620 => x"53442063",
  2621 => x"61726420",
  2622 => x"72657365",
  2623 => x"74206661",
  2624 => x"696c6564",
  2625 => x"210a0000",
  2626 => x"53444843",
  2627 => x"20657272",
  2628 => x"6f72210a",
  2629 => x"00000000",
  2630 => x"57726974",
  2631 => x"65206661",
  2632 => x"696c6564",
  2633 => x"0a000000",
  2634 => x"52656164",
  2635 => x"20666169",
  2636 => x"6c65640a",
  2637 => x"00000000",
  2638 => x"43617264",
  2639 => x"20696e69",
  2640 => x"74206661",
  2641 => x"696c6564",
  2642 => x"0a000000",
  2643 => x"46415431",
  2644 => x"36202020",
  2645 => x"00000000",
  2646 => x"46415433",
  2647 => x"32202020",
  2648 => x"00000000",
  2649 => x"4e6f2070",
  2650 => x"61727469",
  2651 => x"74696f6e",
  2652 => x"20736967",
  2653 => x"0a000000",
  2654 => x"42616420",
  2655 => x"70617274",
  2656 => x"0a000000",
  2657 => x"4261636b",
  2658 => x"00000000",
  2659 => x"00000002",
  2660 => x"00000002",
  2661 => x"0000283c",
  2662 => x"0000035a",
  2663 => x"00000001",
  2664 => x"00002844",
  2665 => x"00000000",
  2666 => x"00000001",
  2667 => x"00002850",
  2668 => x"00000001",
  2669 => x"00000001",
  2670 => x"0000285c",
  2671 => x"00000002",
  2672 => x"00000001",
  2673 => x"00002864",
  2674 => x"00000003",
  2675 => x"00000001",
  2676 => x"00002874",
  2677 => x"00000004",
  2678 => x"00000002",
  2679 => x"00002884",
  2680 => x"0000036e",
  2681 => x"00000002",
  2682 => x"0000288c",
  2683 => x"00000a3f",
  2684 => x"00000002",
  2685 => x"00002894",
  2686 => x"00002800",
  2687 => x"00000002",
  2688 => x"000028a0",
  2689 => x"000014a6",
  2690 => x"00000000",
  2691 => x"00000000",
  2692 => x"00000000",
  2693 => x"00000004",
  2694 => x"000028a8",
  2695 => x"00002a14",
  2696 => x"00000004",
  2697 => x"000028bc",
  2698 => x"00002990",
  2699 => x"00000000",
  2700 => x"00000000",
  2701 => x"00000000",
  2702 => x"00000000",
  2703 => x"00000000",
  2704 => x"00000000",
  2705 => x"00000000",
  2706 => x"00000000",
  2707 => x"00000000",
  2708 => x"00000000",
  2709 => x"00000000",
  2710 => x"00000000",
  2711 => x"00000000",
  2712 => x"00000000",
  2713 => x"00000000",
  2714 => x"00000000",
  2715 => x"00000000",
  2716 => x"00000000",
  2717 => x"00000000",
  2718 => x"00000000",
  2719 => x"00000000",
  2720 => x"00000006",
  2721 => x"00000000",
  2722 => x"00000000",
  2723 => x"00000002",
  2724 => x"00002ef4",
  2725 => x"000025c5",
  2726 => x"00000002",
  2727 => x"00002f12",
  2728 => x"000025c5",
  2729 => x"00000002",
  2730 => x"00002f30",
  2731 => x"000025c5",
  2732 => x"00000002",
  2733 => x"00002f4e",
  2734 => x"000025c5",
  2735 => x"00000002",
  2736 => x"00002f6c",
  2737 => x"000025c5",
  2738 => x"00000002",
  2739 => x"00002f8a",
  2740 => x"000025c5",
  2741 => x"00000002",
  2742 => x"00002fa8",
  2743 => x"000025c5",
  2744 => x"00000002",
  2745 => x"00002fc6",
  2746 => x"000025c5",
  2747 => x"00000002",
  2748 => x"00002fe4",
  2749 => x"000025c5",
  2750 => x"00000002",
  2751 => x"00003002",
  2752 => x"000025c5",
  2753 => x"00000002",
  2754 => x"00003020",
  2755 => x"000025c5",
  2756 => x"00000002",
  2757 => x"0000303e",
  2758 => x"000025c5",
  2759 => x"00000002",
  2760 => x"0000305c",
  2761 => x"000025c5",
  2762 => x"00000004",
  2763 => x"00002984",
  2764 => x"00000000",
  2765 => x"00000000",
  2766 => x"00000000",
  2767 => x"00002785",
  2768 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

