-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity boot_rom is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of boot_rom is


  type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"55",x"AA",x"00",x"00",x"00",x"00",x"1E",x"70", -- 0x0000
    x"00",x"00",x"23",x"80",x"C9",x"00",x"00",x"C9", -- 0x0008
    x"00",x"00",x"C9",x"00",x"00",x"C9",x"00",x"00", -- 0x0010
    x"C9",x"00",x"00",x"C9",x"00",x"00",x"C9",x"00", -- 0x0018
    x"00",x"ED",x"45",x"ED",x"56",x"F3",x"CD",x"41", -- 0x0020
    x"80",x"21",x"33",x"00",x"22",x"C8",x"73",x"CD", -- 0x0028
    x"85",x"1F",x"11",x"00",x"40",x"AF",x"6F",x"67", -- 0x0030
    x"CD",x"82",x"1F",x"CD",x"4A",x"83",x"C3",x"74", -- 0x0038
    x"80",x"21",x"90",x"70",x"11",x"03",x"70",x"CD", -- 0x0040
    x"6A",x"80",x"11",x"00",x"70",x"21",x"0B",x"98", -- 0x0048
    x"01",x"08",x"98",x"CD",x"5F",x"80",x"11",x"90", -- 0x0050
    x"70",x"21",x"AE",x"98",x"01",x"AE",x"98",x"AF", -- 0x0058
    x"ED",x"42",x"C5",x"4D",x"44",x"E1",x"C8",x"ED", -- 0x0060
    x"B0",x"C9",x"AF",x"E5",x"ED",x"52",x"E1",x"C8", -- 0x0068
    x"12",x"13",x"18",x"F7",x"00",x"18",x"FE",x"31", -- 0x0070
    x"8F",x"70",x"CD",x"83",x"80",x"CD",x"4A",x"83", -- 0x0078
    x"C3",x"74",x"80",x"21",x"90",x"70",x"11",x"03", -- 0x0080
    x"70",x"CD",x"AC",x"80",x"11",x"00",x"70",x"21", -- 0x0088
    x"0B",x"98",x"01",x"08",x"98",x"CD",x"A1",x"80", -- 0x0090
    x"11",x"90",x"70",x"21",x"AE",x"98",x"01",x"AE", -- 0x0098
    x"98",x"AF",x"ED",x"42",x"C5",x"4D",x"44",x"E1", -- 0x00A0
    x"C8",x"ED",x"B0",x"C9",x"AF",x"E5",x"ED",x"52", -- 0x00A8
    x"E1",x"C8",x"12",x"13",x"18",x"F7",x"04",x"05", -- 0x00B0
    x"C8",x"CB",x"3A",x"CB",x"1B",x"10",x"FA",x"C9", -- 0x00B8
    x"F5",x"C5",x"E5",x"21",x"00",x"00",x"CB",x"38", -- 0x00C0
    x"CB",x"19",x"38",x"0A",x"78",x"B1",x"28",x"0D", -- 0x00C8
    x"CB",x"23",x"CB",x"12",x"18",x"F0",x"19",x"CB", -- 0x00D0
    x"23",x"CB",x"12",x"18",x"E9",x"EB",x"E1",x"C1", -- 0x00D8
    x"F1",x"C9",x"C5",x"E5",x"F5",x"7C",x"EE",x"80", -- 0x00E0
    x"67",x"78",x"EE",x"80",x"47",x"F1",x"A7",x"ED", -- 0x00E8
    x"42",x"E1",x"C1",x"C9",x"B7",x"C8",x"FE",x"08", -- 0x00F0
    x"38",x"09",x"41",x"4C",x"65",x"2E",x"00",x"D6", -- 0x00F8
    x"08",x"18",x"F2",x"29",x"CB",x"11",x"CB",x"10", -- 0x0100
    x"3D",x"20",x"F8",x"C9",x"B7",x"C8",x"FE",x"08", -- 0x0108
    x"38",x"09",x"6C",x"61",x"48",x"06",x"00",x"D6", -- 0x0110
    x"08",x"18",x"F2",x"CB",x"38",x"CB",x"19",x"CB", -- 0x0118
    x"1C",x"CB",x"1D",x"3D",x"20",x"F5",x"C9",x"E3", -- 0x0120
    x"D5",x"DD",x"E5",x"DD",x"21",x"00",x"00",x"DD", -- 0x0128
    x"39",x"DD",x"56",x"09",x"DD",x"74",x"09",x"DD", -- 0x0130
    x"5E",x"08",x"DD",x"75",x"08",x"D5",x"C5",x"F5", -- 0x0138
    x"21",x"00",x"00",x"11",x"00",x"00",x"06",x"20", -- 0x0140
    x"DD",x"4E",x"FD",x"DD",x"CB",x"FF",x"3E",x"DD", -- 0x0148
    x"CB",x"FE",x"1E",x"DD",x"CB",x"07",x"1E",x"DD", -- 0x0150
    x"CB",x"06",x"1E",x"30",x"12",x"7D",x"DD",x"86", -- 0x0158
    x"04",x"6F",x"7C",x"DD",x"8E",x"05",x"67",x"7B", -- 0x0160
    x"DD",x"8E",x"FC",x"5F",x"7A",x"89",x"57",x"DD", -- 0x0168
    x"CB",x"04",x"26",x"DD",x"CB",x"05",x"16",x"DD", -- 0x0170
    x"CB",x"FC",x"16",x"CB",x"11",x"10",x"CC",x"DD", -- 0x0178
    x"71",x"FD",x"42",x"4B",x"F1",x"D1",x"D1",x"DD", -- 0x0180
    x"E1",x"D1",x"33",x"33",x"33",x"33",x"C9",x"EB", -- 0x0188
    x"E3",x"F5",x"DD",x"E5",x"DD",x"21",x"00",x"00", -- 0x0190
    x"DD",x"39",x"C5",x"D5",x"DD",x"56",x"09",x"DD", -- 0x0198
    x"74",x"09",x"DD",x"5E",x"08",x"DD",x"75",x"08", -- 0x01A0
    x"CD",x"B7",x"81",x"E1",x"C1",x"CD",x"53",x"82", -- 0x01A8
    x"DD",x"E1",x"F1",x"D1",x"33",x"33",x"C9",x"F5", -- 0x01B0
    x"21",x"00",x"00",x"01",x"00",x"00",x"DD",x"36", -- 0x01B8
    x"F8",x"21",x"18",x"02",x"19",x"37",x"DD",x"CB", -- 0x01C0
    x"FC",x"16",x"DD",x"CB",x"FD",x"16",x"DD",x"CB", -- 0x01C8
    x"FE",x"16",x"DD",x"CB",x"FF",x"16",x"DD",x"35", -- 0x01D0
    x"F8",x"28",x"2E",x"CB",x"11",x"CB",x"10",x"CB", -- 0x01D8
    x"15",x"CB",x"14",x"ED",x"52",x"38",x"DD",x"20", -- 0x01E0
    x"10",x"78",x"DD",x"96",x"07",x"38",x"D5",x"20", -- 0x01E8
    x"08",x"79",x"DD",x"96",x"06",x"38",x"CD",x"18", -- 0x01F0
    x"04",x"79",x"DD",x"96",x"06",x"4F",x"78",x"DD", -- 0x01F8
    x"9E",x"07",x"47",x"30",x"C1",x"2B",x"A7",x"18", -- 0x0200
    x"BD",x"F1",x"E5",x"60",x"69",x"C1",x"C9",x"EB", -- 0x0208
    x"E3",x"F5",x"E5",x"21",x"06",x"00",x"39",x"7E", -- 0x0210
    x"A3",x"77",x"23",x"7E",x"A2",x"77",x"D1",x"23", -- 0x0218
    x"7E",x"73",x"A1",x"4F",x"23",x"7E",x"72",x"A0", -- 0x0220
    x"47",x"F1",x"D1",x"E1",x"C9",x"EB",x"E3",x"F5", -- 0x0228
    x"E5",x"21",x"06",x"00",x"39",x"7E",x"B3",x"77", -- 0x0230
    x"23",x"7E",x"B2",x"77",x"D1",x"23",x"7E",x"73", -- 0x0238
    x"B1",x"4F",x"23",x"7E",x"72",x"B0",x"47",x"F1", -- 0x0240
    x"D1",x"E1",x"C9",x"2C",x"C0",x"24",x"C0",x"0C", -- 0x0248
    x"C0",x"04",x"C9",x"F5",x"7D",x"2F",x"6F",x"7C", -- 0x0250
    x"2F",x"67",x"79",x"2F",x"4F",x"78",x"2F",x"47", -- 0x0258
    x"F1",x"C9",x"C5",x"D5",x"5E",x"23",x"56",x"23", -- 0x0260
    x"4E",x"23",x"46",x"EB",x"CD",x"27",x"81",x"C3", -- 0x0268
    x"72",x"82",x"EB",x"70",x"2B",x"71",x"2B",x"72", -- 0x0270
    x"2B",x"73",x"C9",x"F5",x"7E",x"83",x"77",x"5F", -- 0x0278
    x"23",x"7E",x"8A",x"77",x"57",x"23",x"7E",x"89", -- 0x0280
    x"77",x"4F",x"23",x"7E",x"88",x"77",x"47",x"2B", -- 0x0288
    x"2B",x"2B",x"F1",x"C9",x"F5",x"7E",x"93",x"77", -- 0x0290
    x"5F",x"23",x"7E",x"9A",x"77",x"57",x"23",x"7E", -- 0x0298
    x"99",x"77",x"4F",x"23",x"7E",x"98",x"77",x"47", -- 0x02A0
    x"2B",x"2B",x"2B",x"F1",x"C9",x"5E",x"23",x"56", -- 0x02A8
    x"23",x"4E",x"23",x"46",x"EB",x"CD",x"F4",x"80", -- 0x02B0
    x"C3",x"BB",x"82",x"EB",x"70",x"2B",x"71",x"2B", -- 0x02B8
    x"72",x"2B",x"73",x"C9",x"E1",x"C5",x"D5",x"DD", -- 0x02C0
    x"E5",x"DD",x"21",x"00",x"00",x"DD",x"39",x"E9", -- 0x02C8
    x"E1",x"C5",x"D5",x"DD",x"E5",x"DD",x"21",x"00", -- 0x02D0
    x"00",x"DD",x"39",x"5E",x"23",x"56",x"23",x"EB", -- 0x02D8
    x"39",x"F9",x"EB",x"E9",x"DD",x"F9",x"DD",x"E1", -- 0x02E0
    x"D1",x"C1",x"C9",x"DD",x"F9",x"DD",x"E1",x"D1", -- 0x02E8
    x"33",x"33",x"C9",x"F5",x"E5",x"D5",x"C5",x"AF", -- 0x02F0
    x"EB",x"BE",x"ED",x"A0",x"20",x"FB",x"C1",x"D1", -- 0x02F8
    x"E1",x"F1",x"C9",x"E5",x"D5",x"C5",x"F5",x"AF", -- 0x0300
    x"47",x"4F",x"ED",x"B1",x"2B",x"EB",x"BE",x"ED", -- 0x0308
    x"A0",x"20",x"FB",x"F1",x"C1",x"D1",x"E1",x"C9", -- 0x0310
    x"7E",x"BB",x"C8",x"B7",x"23",x"20",x"F9",x"21", -- 0x0318
    x"00",x"00",x"C9",x"CD",x"D0",x"82",x"00",x"00", -- 0x0320
    x"21",x"0B",x"98",x"E5",x"0E",x"12",x"1E",x"0C", -- 0x0328
    x"CD",x"64",x"97",x"E1",x"11",x"00",x"00",x"01", -- 0x0330
    x"50",x"C3",x"6B",x"62",x"A7",x"ED",x"42",x"30", -- 0x0338
    x"03",x"13",x"18",x"F3",x"C3",x"00",x"00",x"C3", -- 0x0340
    x"E4",x"82",x"CD",x"D0",x"82",x"A0",x"FF",x"FD", -- 0x0348
    x"E5",x"CD",x"00",x"98",x"CD",x"F8",x"97",x"CD", -- 0x0350
    x"2C",x"89",x"1E",x"00",x"CD",x"01",x"86",x"1E", -- 0x0358
    x"F4",x"CD",x"E6",x"97",x"CD",x"13",x"86",x"CD", -- 0x0360
    x"D6",x"97",x"3E",x"0B",x"01",x"24",x"00",x"ED", -- 0x0368
    x"79",x"21",x"3E",x"00",x"39",x"EB",x"CD",x"1E", -- 0x0370
    x"8F",x"B7",x"28",x"04",x"5F",x"CD",x"23",x"83", -- 0x0378
    x"11",x"1C",x"98",x"CD",x"5E",x"92",x"B7",x"28", -- 0x0380
    x"04",x"5F",x"CD",x"23",x"83",x"DD",x"70",x"A2", -- 0x0388
    x"CD",x"F1",x"85",x"21",x"25",x"98",x"E5",x"0E", -- 0x0390
    x"01",x"1E",x"03",x"CD",x"64",x"97",x"E1",x"21", -- 0x0398
    x"41",x"98",x"E5",x"0E",x"03",x"59",x"CD",x"64", -- 0x03A0
    x"97",x"E1",x"21",x"5A",x"98",x"E5",x"0E",x"14", -- 0x03A8
    x"1E",x"01",x"CD",x"64",x"97",x"E1",x"21",x"78", -- 0x03B0
    x"98",x"E5",x"0E",x"16",x"1E",x"01",x"CD",x"64", -- 0x03B8
    x"97",x"E1",x"DD",x"36",x"A3",x"00",x"21",x"0C", -- 0x03C0
    x"00",x"39",x"E5",x"01",x"1B",x"00",x"11",x"03", -- 0x03C8
    x"70",x"CD",x"02",x"93",x"E1",x"B7",x"20",x"2C", -- 0x03D0
    x"DD",x"7E",x"AA",x"DD",x"B6",x"AB",x"28",x"24", -- 0x03D8
    x"DD",x"34",x"A3",x"11",x"3B",x"00",x"21",x"03", -- 0x03E0
    x"70",x"CD",x"18",x"83",x"72",x"21",x"03",x"70", -- 0x03E8
    x"E5",x"DD",x"7E",x"A3",x"C6",x"04",x"4F",x"1E", -- 0x03F0
    x"04",x"CD",x"64",x"97",x"E1",x"DD",x"7E",x"A3", -- 0x03F8
    x"FE",x"0A",x"20",x"C2",x"21",x"00",x"70",x"E5", -- 0x0400
    x"0E",x"05",x"CD",x"E3",x"85",x"E1",x"DD",x"36", -- 0x0408
    x"A1",x"05",x"DD",x"36",x"A4",x"00",x"1E",x"00", -- 0x0410
    x"CD",x"B7",x"97",x"DD",x"75",x"A6",x"DD",x"74", -- 0x0418
    x"A7",x"CB",x"55",x"28",x"2D",x"DD",x"4E",x"A3", -- 0x0420
    x"06",x"00",x"21",x"04",x"00",x"09",x"4D",x"44", -- 0x0428
    x"DD",x"6E",x"A1",x"26",x"00",x"CD",x"E2",x"80", -- 0x0430
    x"30",x"18",x"21",x"96",x"98",x"E5",x"CD",x"E0", -- 0x0438
    x"85",x"E1",x"DD",x"34",x"A1",x"21",x"00",x"70", -- 0x0440
    x"E5",x"CD",x"E0",x"85",x"E1",x"DD",x"34",x"A4", -- 0x0448
    x"18",x"58",x"DD",x"CB",x"A6",x"46",x"28",x"1F", -- 0x0450
    x"3E",x"05",x"DD",x"BE",x"A1",x"30",x"18",x"21", -- 0x0458
    x"96",x"98",x"E5",x"CD",x"E0",x"85",x"E1",x"DD", -- 0x0460
    x"35",x"A1",x"21",x"00",x"70",x"E5",x"CD",x"E0", -- 0x0468
    x"85",x"E1",x"DD",x"35",x"A4",x"18",x"33",x"DD", -- 0x0470
    x"CB",x"A6",x"5E",x"28",x"0B",x"AF",x"DD",x"B6", -- 0x0478
    x"A2",x"28",x"0E",x"DD",x"35",x"A2",x"18",x"09", -- 0x0480
    x"DD",x"CB",x"A6",x"4E",x"28",x"1C",x"DD",x"34", -- 0x0488
    x"A2",x"DD",x"4E",x"A2",x"06",x"00",x"11",x"0E", -- 0x0490
    x"01",x"CD",x"C0",x"80",x"7A",x"07",x"9F",x"4F", -- 0x0498
    x"41",x"CD",x"EF",x"94",x"DD",x"36",x"A5",x"00", -- 0x04A0
    x"18",x"34",x"DD",x"7E",x"A7",x"2E",x"00",x"E6", -- 0x04A8
    x"C0",x"67",x"7D",x"B4",x"28",x"06",x"DD",x"36", -- 0x04B0
    x"A5",x"01",x"18",x"22",x"AF",x"DD",x"77",x"AC", -- 0x04B8
    x"DD",x"77",x"AD",x"01",x"F0",x"0A",x"DD",x"6E", -- 0x04C0
    x"AC",x"DD",x"66",x"AD",x"A7",x"ED",x"42",x"30", -- 0x04C8
    x"0A",x"DD",x"34",x"AC",x"20",x"ED",x"DD",x"34", -- 0x04D0
    x"AD",x"18",x"E8",x"C3",x"16",x"84",x"AF",x"DD", -- 0x04D8
    x"B6",x"A5",x"CA",x"90",x"83",x"3E",x"80",x"DD", -- 0x04E0
    x"AE",x"A7",x"DD",x"B6",x"A6",x"CA",x"B7",x"85", -- 0x04E8
    x"DD",x"4E",x"A4",x"06",x"00",x"11",x"1B",x"00", -- 0x04F0
    x"CD",x"C0",x"80",x"D5",x"DD",x"4E",x"A2",x"11", -- 0x04F8
    x"0E",x"01",x"CD",x"C0",x"80",x"EB",x"D1",x"19", -- 0x0500
    x"0E",x"11",x"09",x"EB",x"7A",x"07",x"9F",x"4F", -- 0x0508
    x"41",x"CD",x"EF",x"94",x"21",x"0C",x"00",x"39", -- 0x0510
    x"E5",x"01",x"0D",x"00",x"11",x"03",x"70",x"CD", -- 0x0518
    x"02",x"93",x"E1",x"11",x"0D",x"00",x"21",x"03", -- 0x0520
    x"70",x"CD",x"18",x"83",x"7D",x"B4",x"28",x"01", -- 0x0528
    x"72",x"1E",x"20",x"21",x"03",x"70",x"CD",x"18", -- 0x0530
    x"83",x"7D",x"B4",x"28",x"01",x"72",x"11",x"03", -- 0x0538
    x"70",x"21",x"14",x"00",x"39",x"CD",x"F3",x"82", -- 0x0540
    x"11",x"99",x"98",x"21",x"14",x"00",x"39",x"CD", -- 0x0548
    x"03",x"83",x"21",x"9E",x"98",x"E5",x"0E",x"12", -- 0x0550
    x"1E",x"04",x"CD",x"64",x"97",x"E1",x"21",x"14", -- 0x0558
    x"00",x"39",x"E5",x"0E",x"12",x"1E",x"0C",x"CD", -- 0x0560
    x"64",x"97",x"E1",x"11",x"A6",x"98",x"21",x"24", -- 0x0568
    x"00",x"39",x"CD",x"F3",x"82",x"21",x"14",x"00", -- 0x0570
    x"39",x"EB",x"21",x"24",x"00",x"39",x"CD",x"03", -- 0x0578
    x"83",x"EB",x"CD",x"5E",x"92",x"B7",x"28",x"04", -- 0x0580
    x"5F",x"CD",x"23",x"83",x"FD",x"21",x"00",x"80", -- 0x0588
    x"21",x"0C",x"00",x"39",x"E5",x"01",x"00",x"80", -- 0x0590
    x"FD",x"E5",x"D1",x"CD",x"02",x"93",x"E1",x"DD", -- 0x0598
    x"77",x"A0",x"B7",x"20",x"08",x"DD",x"7E",x"AA", -- 0x05A0
    x"DD",x"B6",x"AB",x"20",x"E3",x"AF",x"DD",x"B6", -- 0x05A8
    x"A0",x"28",x"04",x"5F",x"CD",x"23",x"83",x"FD", -- 0x05B0
    x"21",x"01",x"71",x"3E",x"3E",x"32",x"00",x"71", -- 0x05B8
    x"FD",x"36",x"00",x"04",x"FD",x"36",x"01",x"D3", -- 0x05C0
    x"FD",x"36",x"02",x"24",x"FD",x"36",x"03",x"C3", -- 0x05C8
    x"FD",x"36",x"04",x"00",x"FD",x"36",x"05",x"00", -- 0x05D0
    x"C3",x"00",x"71",x"FD",x"E1",x"C3",x"E4",x"82", -- 0x05D8
    x"DD",x"4E",x"A1",x"1E",x"02",x"C3",x"64",x"97", -- 0x05E0
    x"CD",x"C0",x"08",x"2A",x"F6",x"73",x"19",x"EB", -- 0x05E8
    x"C9",x"DD",x"E5",x"2A",x"F6",x"73",x"11",x"00", -- 0x05F0
    x"03",x"3E",x"20",x"CD",x"82",x"1F",x"DD",x"E1", -- 0x05F8
    x"C9",x"CD",x"C4",x"82",x"DD",x"7E",x"02",x"21", -- 0x0600
    x"00",x"00",x"11",x"00",x"40",x"CD",x"82",x"1F", -- 0x0608
    x"C3",x"E4",x"82",x"DD",x"E5",x"CD",x"7F",x"1F", -- 0x0610
    x"DD",x"E1",x"C9",x"CD",x"D0",x"82",x"00",x"00", -- 0x0618
    x"11",x"00",x"00",x"DD",x"4E",x"02",x"DD",x"46", -- 0x0620
    x"03",x"6B",x"62",x"A7",x"ED",x"42",x"30",x"03", -- 0x0628
    x"13",x"18",x"F0",x"C3",x"E4",x"82",x"CD",x"C4", -- 0x0630
    x"82",x"01",x"51",x"00",x"ED",x"59",x"C3",x"E4", -- 0x0638
    x"82",x"C5",x"D5",x"3E",x"FF",x"01",x"51",x"00", -- 0x0640
    x"ED",x"79",x"0B",x"ED",x"50",x"7A",x"D1",x"C1", -- 0x0648
    x"C9",x"C5",x"DD",x"E5",x"D5",x"DD",x"E1",x"3E", -- 0x0650
    x"FF",x"01",x"51",x"00",x"ED",x"79",x"DD",x"2B", -- 0x0658
    x"DD",x"E5",x"E1",x"7D",x"B4",x"20",x"F0",x"DD", -- 0x0660
    x"E1",x"C1",x"C9",x"C5",x"CD",x"71",x"86",x"C1", -- 0x0668
    x"C9",x"3E",x"01",x"01",x"50",x"00",x"ED",x"79", -- 0x0670
    x"C3",x"41",x"86",x"CD",x"D0",x"82",x"FE",x"FF", -- 0x0678
    x"DD",x"CB",x"02",x"7E",x"28",x"19",x"DD",x"CB", -- 0x0680
    x"02",x"BE",x"21",x"00",x"00",x"E5",x"E5",x"1E", -- 0x0688
    x"77",x"CD",x"7B",x"86",x"E1",x"E1",x"DD",x"77", -- 0x0690
    x"FF",x"47",x"3E",x"01",x"B8",x"38",x"5B",x"CD", -- 0x0698
    x"71",x"86",x"AF",x"CD",x"76",x"86",x"DD",x"5E", -- 0x06A0
    x"02",x"CD",x"36",x"86",x"DD",x"4E",x"0A",x"DD", -- 0x06A8
    x"5E",x"0B",x"CD",x"36",x"86",x"59",x"CD",x"36", -- 0x06B0
    x"86",x"DD",x"5E",x"09",x"CD",x"36",x"86",x"DD", -- 0x06B8
    x"5E",x"08",x"CD",x"36",x"86",x"DD",x"36",x"FE", -- 0x06C0
    x"01",x"DD",x"7E",x"02",x"FE",x"40",x"20",x"04", -- 0x06C8
    x"DD",x"36",x"FE",x"95",x"FE",x"48",x"20",x"04", -- 0x06D0
    x"DD",x"36",x"FE",x"87",x"DD",x"5E",x"FE",x"CD", -- 0x06D8
    x"36",x"86",x"DD",x"36",x"FE",x"0A",x"CD",x"41", -- 0x06E0
    x"86",x"DD",x"77",x"FF",x"B7",x"F2",x"FA",x"86", -- 0x06E8
    x"DD",x"35",x"FE",x"DD",x"46",x"FE",x"04",x"05", -- 0x06F0
    x"20",x"EC",x"DD",x"7E",x"FF",x"C3",x"E4",x"82", -- 0x06F8
    x"CD",x"D0",x"82",x"F6",x"FF",x"3E",x"01",x"01", -- 0x0700
    x"50",x"00",x"ED",x"79",x"11",x"64",x"00",x"CD", -- 0x0708
    x"51",x"86",x"DD",x"70",x"F7",x"68",x"60",x"E5", -- 0x0710
    x"E5",x"1E",x"40",x"CD",x"7B",x"86",x"E1",x"E1", -- 0x0718
    x"3D",x"C2",x"25",x"88",x"68",x"60",x"E5",x"21", -- 0x0720
    x"AA",x"01",x"E5",x"1E",x"48",x"CD",x"7B",x"86", -- 0x0728
    x"E1",x"E1",x"3D",x"C2",x"CA",x"87",x"DD",x"70", -- 0x0730
    x"F6",x"DD",x"7E",x"F6",x"FE",x"04",x"30",x"11", -- 0x0738
    x"4F",x"21",x"04",x"00",x"39",x"09",x"E5",x"CD", -- 0x0740
    x"41",x"86",x"E1",x"77",x"DD",x"34",x"F6",x"18", -- 0x0748
    x"E8",x"DD",x"46",x"FC",x"05",x"C2",x"25",x"88", -- 0x0750
    x"DD",x"7E",x"FD",x"FE",x"AA",x"C2",x"25",x"88", -- 0x0758
    x"DD",x"36",x"F8",x"E8",x"DD",x"36",x"F9",x"03", -- 0x0760
    x"DD",x"7E",x"F8",x"DD",x"B6",x"F9",x"28",x"15", -- 0x0768
    x"21",x"00",x"40",x"E5",x"65",x"E5",x"1E",x"E9", -- 0x0770
    x"CD",x"7B",x"86",x"E1",x"E1",x"B7",x"28",x"05", -- 0x0778
    x"CD",x"3B",x"88",x"18",x"E3",x"DD",x"7E",x"F8", -- 0x0780
    x"DD",x"B6",x"F9",x"28",x"3B",x"21",x"00",x"00", -- 0x0788
    x"E5",x"E5",x"1E",x"7A",x"CD",x"7B",x"86",x"E1", -- 0x0790
    x"E1",x"B7",x"20",x"2C",x"DD",x"77",x"F6",x"DD", -- 0x0798
    x"7E",x"F6",x"FE",x"04",x"30",x"13",x"4F",x"06", -- 0x07A0
    x"00",x"21",x"04",x"00",x"39",x"09",x"E5",x"CD", -- 0x07A8
    x"41",x"86",x"E1",x"77",x"DD",x"34",x"F6",x"18", -- 0x07B0
    x"E6",x"DD",x"CB",x"FA",x"76",x"28",x"04",x"3E", -- 0x07B8
    x"0C",x"18",x"02",x"3E",x"04",x"DD",x"77",x"F7", -- 0x07C0
    x"18",x"5B",x"68",x"60",x"E5",x"E5",x"1E",x"E9", -- 0x07C8
    x"CD",x"7B",x"86",x"E1",x"E1",x"47",x"3E",x"01", -- 0x07D0
    x"B8",x"38",x"06",x"DD",x"36",x"F7",x"02",x"18", -- 0x07D8
    x"03",x"DD",x"77",x"F7",x"DD",x"36",x"F8",x"E8", -- 0x07E0
    x"DD",x"36",x"F9",x"03",x"DD",x"7E",x"F8",x"DD", -- 0x07E8
    x"B6",x"F9",x"28",x"14",x"21",x"00",x"00",x"E5", -- 0x07F0
    x"E5",x"1E",x"E9",x"CD",x"7B",x"86",x"E1",x"E1", -- 0x07F8
    x"B7",x"28",x"05",x"CD",x"3B",x"88",x"18",x"E4", -- 0x0800
    x"DD",x"7E",x"F8",x"DD",x"B6",x"F9",x"28",x"11", -- 0x0808
    x"21",x"00",x"00",x"E5",x"26",x"02",x"E5",x"1E", -- 0x0810
    x"50",x"CD",x"7B",x"86",x"E1",x"E1",x"B7",x"28", -- 0x0818
    x"04",x"DD",x"36",x"F7",x"00",x"DD",x"46",x"F7", -- 0x0820
    x"78",x"32",x"8D",x"70",x"CD",x"6B",x"86",x"04", -- 0x0828
    x"05",x"28",x"03",x"AF",x"18",x"02",x"3E",x"01", -- 0x0830
    x"C3",x"E4",x"82",x"11",x"E8",x"03",x"CD",x"1B", -- 0x0838
    x"86",x"DD",x"6E",x"F8",x"DD",x"66",x"F9",x"2B", -- 0x0840
    x"DD",x"75",x"F8",x"DD",x"74",x"F9",x"C9",x"CD", -- 0x0848
    x"D0",x"82",x"FC",x"FF",x"FD",x"E5",x"DD",x"5E", -- 0x0850
    x"0E",x"DD",x"56",x"0F",x"3A",x"8D",x"70",x"CB", -- 0x0858
    x"5F",x"20",x"0B",x"D5",x"21",x"10",x"00",x"39", -- 0x0860
    x"3E",x"09",x"CD",x"AD",x"82",x"D1",x"DD",x"36", -- 0x0868
    x"FD",x"01",x"D5",x"DD",x"6E",x"0A",x"DD",x"66", -- 0x0870
    x"0B",x"E5",x"DD",x"6E",x"08",x"DD",x"66",x"09", -- 0x0878
    x"E5",x"1E",x"51",x"CD",x"7B",x"86",x"E1",x"E1", -- 0x0880
    x"B7",x"D1",x"C2",x"0E",x"89",x"FD",x"21",x"E8", -- 0x0888
    x"03",x"D5",x"11",x"64",x"00",x"CD",x"1B",x"86", -- 0x0890
    x"D1",x"CD",x"41",x"86",x"DD",x"77",x"FC",x"3C", -- 0x0898
    x"20",x"09",x"FD",x"2B",x"FD",x"E5",x"E1",x"7D", -- 0x08A0
    x"B4",x"20",x"E6",x"DD",x"46",x"FC",x"04",x"04", -- 0x08A8
    x"20",x"5C",x"DD",x"4E",x"0C",x"DD",x"46",x"0D", -- 0x08B0
    x"21",x"02",x"02",x"A7",x"ED",x"42",x"A7",x"ED", -- 0x08B8
    x"52",x"DD",x"75",x"FE",x"DD",x"74",x"FF",x"79", -- 0x08C0
    x"B0",x"28",x"0B",x"D5",x"DD",x"5E",x"0C",x"DD", -- 0x08C8
    x"56",x"0D",x"CD",x"51",x"86",x"D1",x"DD",x"7E", -- 0x08D0
    x"02",x"DD",x"B6",x"03",x"28",x"1B",x"DD",x"6E", -- 0x08D8
    x"02",x"DD",x"66",x"03",x"23",x"DD",x"75",x"02", -- 0x08E0
    x"DD",x"74",x"03",x"2B",x"E5",x"CD",x"41",x"86", -- 0x08E8
    x"E1",x"77",x"1B",x"7B",x"B2",x"20",x"E7",x"18", -- 0x08F0
    x"08",x"CD",x"41",x"86",x"1B",x"7B",x"B2",x"20", -- 0x08F8
    x"F8",x"DD",x"5E",x"FE",x"DD",x"56",x"FF",x"CD", -- 0x0900
    x"51",x"86",x"DD",x"36",x"FD",x"00",x"CD",x"6B", -- 0x0908
    x"86",x"DD",x"7E",x"FD",x"FD",x"E1",x"C3",x"E4", -- 0x0910
    x"82",x"DD",x"E5",x"3A",x"C4",x"73",x"F6",x"20", -- 0x0918
    x"4F",x"06",x"01",x"CD",x"D9",x"1F",x"CD",x"DC", -- 0x0920
    x"1F",x"DD",x"E1",x"C9",x"DD",x"E5",x"3A",x"C4", -- 0x0928
    x"73",x"E6",x"DF",x"4F",x"06",x"01",x"CD",x"D9", -- 0x0930
    x"1F",x"DD",x"E1",x"C9",x"CD",x"D0",x"82",x"00", -- 0x0938
    x"00",x"FD",x"E5",x"DD",x"5E",x"08",x"DD",x"56", -- 0x0940
    x"09",x"DD",x"6E",x"02",x"DD",x"66",x"03",x"E5", -- 0x0948
    x"FD",x"E1",x"7B",x"62",x"1B",x"B4",x"28",x"0A", -- 0x0950
    x"DD",x"46",x"04",x"FD",x"70",x"00",x"FD",x"23", -- 0x0958
    x"18",x"F0",x"FD",x"E1",x"C3",x"E4",x"82",x"CD", -- 0x0960
    x"D0",x"82",x"FE",x"FF",x"FD",x"E5",x"DD",x"6E", -- 0x0968
    x"02",x"DD",x"66",x"03",x"E5",x"FD",x"E1",x"59", -- 0x0970
    x"50",x"AF",x"DD",x"77",x"FE",x"DD",x"77",x"FF", -- 0x0978
    x"DD",x"6E",x"08",x"DD",x"66",x"09",x"2B",x"DD", -- 0x0980
    x"75",x"08",x"DD",x"74",x"09",x"23",x"7D",x"B4", -- 0x0988
    x"28",x"18",x"6B",x"62",x"13",x"4E",x"06",x"00", -- 0x0990
    x"60",x"FD",x"6E",x"00",x"ED",x"42",x"DD",x"75", -- 0x0998
    x"FE",x"DD",x"74",x"FF",x"7D",x"B4",x"FD",x"23", -- 0x09A0
    x"28",x"D6",x"DD",x"6E",x"FE",x"DD",x"66",x"FF", -- 0x09A8
    x"FD",x"E1",x"C3",x"E4",x"82",x"CD",x"D0",x"82", -- 0x09B0
    x"FC",x"FF",x"FD",x"E5",x"FD",x"2A",x"8E",x"70", -- 0x09B8
    x"01",x"02",x"00",x"DD",x"6E",x"02",x"DD",x"66", -- 0x09C0
    x"03",x"A7",x"ED",x"42",x"38",x"56",x"FD",x"4E", -- 0x09C8
    x"06",x"FD",x"46",x"07",x"DD",x"6E",x"02",x"DD", -- 0x09D0
    x"66",x"03",x"ED",x"42",x"30",x"46",x"FD",x"7E", -- 0x09D8
    x"00",x"FE",x"02",x"20",x"3F",x"21",x"02",x"00", -- 0x09E0
    x"E5",x"DD",x"6E",x"02",x"29",x"E5",x"FD",x"6E", -- 0x09E8
    x"0A",x"FD",x"66",x"0B",x"E5",x"FD",x"6E",x"08", -- 0x09F0
    x"FD",x"66",x"09",x"E5",x"DD",x"6E",x"03",x"26", -- 0x09F8
    x"00",x"5C",x"54",x"C1",x"09",x"EB",x"C1",x"ED", -- 0x0A00
    x"4A",x"E5",x"D5",x"21",x"0A",x"00",x"39",x"EB", -- 0x0A08
    x"CD",x"4F",x"88",x"E1",x"E1",x"E1",x"E1",x"B7", -- 0x0A10
    x"20",x"0A",x"DD",x"66",x"FD",x"DD",x"5E",x"FC", -- 0x0A18
    x"B3",x"6F",x"18",x"03",x"21",x"01",x"00",x"FD", -- 0x0A20
    x"E1",x"C3",x"E4",x"82",x"FD",x"E5",x"DD",x"E5", -- 0x0A28
    x"D5",x"FD",x"E1",x"DD",x"2A",x"8E",x"70",x"21", -- 0x0A30
    x"06",x"00",x"ED",x"4B",x"8E",x"70",x"09",x"46", -- 0x0A38
    x"23",x"66",x"68",x"01",x"FE",x"FF",x"09",x"4D", -- 0x0A40
    x"44",x"FD",x"2B",x"FD",x"2B",x"FD",x"E5",x"E1", -- 0x0A48
    x"A7",x"ED",x"42",x"38",x"07",x"01",x"00",x"00", -- 0x0A50
    x"69",x"60",x"18",x"26",x"DD",x"6E",x"02",x"01", -- 0x0A58
    x"00",x"00",x"61",x"C5",x"E5",x"FD",x"E5",x"E1", -- 0x0A60
    x"CD",x"27",x"81",x"C5",x"E5",x"DD",x"6E",x"10", -- 0x0A68
    x"DD",x"66",x"11",x"C1",x"09",x"EB",x"DD",x"6E", -- 0x0A70
    x"12",x"DD",x"66",x"13",x"C1",x"ED",x"4A",x"4D", -- 0x0A78
    x"44",x"EB",x"DD",x"E1",x"FD",x"E1",x"C9",x"C5", -- 0x0A80
    x"FD",x"E5",x"DD",x"E5",x"F5",x"D5",x"FD",x"E1", -- 0x0A88
    x"DD",x"2A",x"8E",x"70",x"EB",x"AF",x"77",x"23", -- 0x0A90
    x"77",x"6F",x"67",x"39",x"FD",x"4E",x"04",x"71", -- 0x0A98
    x"FD",x"46",x"05",x"23",x"70",x"3E",x"01",x"A9", -- 0x0AA0
    x"B0",x"28",x"0F",x"DD",x"4E",x"06",x"DD",x"46", -- 0x0AA8
    x"07",x"2B",x"56",x"23",x"66",x"6A",x"ED",x"42", -- 0x0AB0
    x"38",x"04",x"3E",x"01",x"18",x"54",x"AF",x"28", -- 0x0AB8
    x"19",x"6F",x"67",x"39",x"7A",x"23",x"B6",x"20", -- 0x0AC0
    x"11",x"DD",x"7E",x"00",x"FE",x"03",x"20",x"0A", -- 0x0AC8
    x"2B",x"DD",x"4E",x"0C",x"71",x"DD",x"46",x"0D", -- 0x0AD0
    x"23",x"70",x"21",x"00",x"00",x"39",x"46",x"FD", -- 0x0AD8
    x"70",x"06",x"23",x"66",x"FD",x"74",x"07",x"21", -- 0x0AE0
    x"00",x"00",x"39",x"78",x"23",x"B6",x"28",x"09", -- 0x0AE8
    x"2B",x"58",x"23",x"56",x"CD",x"2C",x"8A",x"18", -- 0x0AF0
    x"0C",x"DD",x"4E",x"0E",x"DD",x"46",x"0F",x"DD", -- 0x0AF8
    x"6E",x"0C",x"DD",x"66",x"0D",x"FD",x"75",x"08", -- 0x0B00
    x"FD",x"74",x"09",x"FD",x"71",x"0A",x"FD",x"70", -- 0x0B08
    x"0B",x"AF",x"E1",x"DD",x"E1",x"FD",x"E1",x"C1", -- 0x0B10
    x"C9",x"C5",x"FD",x"E5",x"DD",x"E5",x"F5",x"F5", -- 0x0B18
    x"D5",x"DD",x"E1",x"FD",x"2A",x"8E",x"70",x"21", -- 0x0B20
    x"00",x"00",x"39",x"1A",x"4F",x"13",x"1A",x"47", -- 0x0B28
    x"03",x"71",x"23",x"70",x"79",x"B0",x"28",x"49", -- 0x0B30
    x"DD",x"7E",x"08",x"DD",x"B6",x"09",x"DD",x"B6", -- 0x0B38
    x"0A",x"DD",x"B6",x"0B",x"28",x"3B",x"79",x"E6", -- 0x0B40
    x"0F",x"C2",x"F7",x"8B",x"DD",x"6E",x"08",x"DD", -- 0x0B48
    x"66",x"09",x"DD",x"4E",x"0A",x"DD",x"46",x"0B", -- 0x0B50
    x"CD",x"4B",x"82",x"DD",x"75",x"08",x"DD",x"74", -- 0x0B58
    x"09",x"DD",x"71",x"0A",x"DD",x"70",x"0B",x"DD", -- 0x0B60
    x"7E",x"06",x"DD",x"B6",x"07",x"20",x"14",x"FD", -- 0x0B68
    x"4E",x"04",x"FD",x"46",x"05",x"6F",x"67",x"39", -- 0x0B70
    x"56",x"23",x"66",x"6A",x"A7",x"ED",x"42",x"38", -- 0x0B78
    x"76",x"18",x"4D",x"06",x"04",x"21",x"00",x"00", -- 0x0B80
    x"39",x"5E",x"23",x"56",x"CD",x"B6",x"80",x"FD", -- 0x0B88
    x"4E",x"02",x"06",x"00",x"0B",x"7B",x"A1",x"67", -- 0x0B90
    x"7A",x"A0",x"B4",x"20",x"5A",x"21",x"02",x"00", -- 0x0B98
    x"39",x"E5",x"DD",x"5E",x"06",x"DD",x"56",x"07", -- 0x0BA0
    x"CD",x"B5",x"89",x"4D",x"44",x"E1",x"71",x"23", -- 0x0BA8
    x"70",x"21",x"01",x"00",x"A7",x"ED",x"42",x"38", -- 0x0BB0
    x"04",x"3E",x"01",x"18",x"4B",x"FD",x"4E",x"06", -- 0x0BB8
    x"FD",x"46",x"07",x"21",x"02",x"00",x"39",x"56", -- 0x0BC0
    x"23",x"66",x"6A",x"A7",x"ED",x"42",x"38",x"04", -- 0x0BC8
    x"3E",x"03",x"18",x"34",x"21",x"02",x"00",x"39", -- 0x0BD0
    x"42",x"DD",x"70",x"06",x"23",x"66",x"DD",x"74", -- 0x0BD8
    x"07",x"21",x"02",x"00",x"39",x"58",x"23",x"56", -- 0x0BE0
    x"CD",x"2C",x"8A",x"DD",x"75",x"08",x"DD",x"74", -- 0x0BE8
    x"09",x"DD",x"71",x"0A",x"DD",x"70",x"0B",x"21", -- 0x0BF0
    x"00",x"00",x"39",x"46",x"23",x"66",x"68",x"E5", -- 0x0BF8
    x"DD",x"E5",x"E1",x"C1",x"71",x"23",x"70",x"AF", -- 0x0C00
    x"E1",x"E1",x"DD",x"E1",x"FD",x"E1",x"C1",x"C9", -- 0x0C08
    x"FD",x"E5",x"DD",x"E5",x"F5",x"D5",x"DD",x"E1", -- 0x0C10
    x"C5",x"FD",x"E1",x"CD",x"87",x"8A",x"21",x"00", -- 0x0C18
    x"00",x"39",x"77",x"AF",x"B6",x"20",x"6A",x"21", -- 0x0C20
    x"20",x"00",x"E5",x"DD",x"7E",x"00",x"E6",x"0F", -- 0x0C28
    x"6F",x"29",x"29",x"29",x"29",x"29",x"E5",x"DD", -- 0x0C30
    x"6E",x"0A",x"DD",x"66",x"0B",x"E5",x"DD",x"6E", -- 0x0C38
    x"08",x"DD",x"66",x"09",x"E5",x"FD",x"E5",x"D1", -- 0x0C40
    x"CD",x"4F",x"88",x"E1",x"E1",x"E1",x"E1",x"B7", -- 0x0C48
    x"28",x"02",x"3E",x"01",x"21",x"00",x"00",x"39", -- 0x0C50
    x"77",x"AF",x"B6",x"20",x"34",x"FD",x"46",x"00", -- 0x0C58
    x"B0",x"20",x"04",x"36",x"03",x"18",x"2A",x"FD", -- 0x0C60
    x"CB",x"0B",x"5E",x"20",x"15",x"21",x"0B",x"00", -- 0x0C68
    x"E5",x"DD",x"4E",x"02",x"DD",x"46",x"03",x"FD", -- 0x0C70
    x"E5",x"D1",x"CD",x"67",x"89",x"F1",x"7D",x"B4", -- 0x0C78
    x"28",x"0F",x"DD",x"E5",x"D1",x"CD",x"19",x"8B", -- 0x0C80
    x"21",x"00",x"00",x"39",x"77",x"AF",x"B6",x"28", -- 0x0C88
    x"96",x"21",x"00",x"00",x"39",x"7E",x"E1",x"DD", -- 0x0C90
    x"E1",x"FD",x"E1",x"C9",x"CD",x"D0",x"82",x"FA", -- 0x0C98
    x"FF",x"FD",x"E5",x"DD",x"6E",x"02",x"DD",x"66", -- 0x0CA0
    x"03",x"23",x"23",x"7E",x"23",x"66",x"6F",x"E5", -- 0x0CA8
    x"FD",x"E1",x"01",x"0B",x"00",x"C5",x"0E",x"20", -- 0x0CB0
    x"EB",x"CD",x"3C",x"89",x"E1",x"DD",x"6E",x"04", -- 0x0CB8
    x"DD",x"66",x"05",x"46",x"23",x"66",x"68",x"EB", -- 0x0CC0
    x"DD",x"36",x"FB",x"00",x"DD",x"36",x"FC",x"00", -- 0x0CC8
    x"DD",x"36",x"FD",x"08",x"DD",x"4E",x"FC",x"DD", -- 0x0CD0
    x"34",x"FC",x"06",x"00",x"6B",x"62",x"09",x"46", -- 0x0CD8
    x"DD",x"70",x"FA",x"3E",x"20",x"B8",x"30",x"05", -- 0x0CE0
    x"78",x"FE",x"2F",x"20",x"03",x"C3",x"79",x"8D", -- 0x0CE8
    x"FE",x"2E",x"28",x"08",x"DD",x"7E",x"FB",x"DD", -- 0x0CF0
    x"BE",x"FD",x"38",x"16",x"DD",x"7E",x"FD",x"FE", -- 0x0CF8
    x"08",x"20",x"76",x"78",x"FE",x"2E",x"20",x"71", -- 0x0D00
    x"DD",x"36",x"FB",x"08",x"DD",x"36",x"FD",x"0B", -- 0x0D08
    x"18",x"C2",x"AF",x"28",x"3B",x"DD",x"4E",x"FD", -- 0x0D10
    x"47",x"0B",x"DD",x"6E",x"FB",x"67",x"CD",x"E2", -- 0x0D18
    x"80",x"30",x"2D",x"DD",x"4E",x"FC",x"DD",x"34", -- 0x0D20
    x"FC",x"44",x"6B",x"62",x"09",x"46",x"DD",x"70", -- 0x0D28
    x"FE",x"DD",x"4E",x"FB",x"DD",x"34",x"FB",x"47", -- 0x0D30
    x"FD",x"E5",x"E1",x"09",x"DD",x"46",x"FA",x"70", -- 0x0D38
    x"DD",x"4E",x"FB",x"DD",x"34",x"FB",x"47",x"FD", -- 0x0D40
    x"E5",x"E1",x"09",x"DD",x"46",x"FE",x"18",x"25", -- 0x0D48
    x"DD",x"7E",x"FA",x"FE",x"61",x"38",x"0F",x"3E", -- 0x0D50
    x"7A",x"DD",x"BE",x"FA",x"38",x"08",x"21",x"02", -- 0x0D58
    x"00",x"39",x"7E",x"D6",x"20",x"77",x"DD",x"4E", -- 0x0D60
    x"FB",x"DD",x"34",x"FB",x"06",x"00",x"FD",x"E5", -- 0x0D68
    x"E1",x"09",x"DD",x"46",x"FA",x"70",x"C3",x"D4", -- 0x0D70
    x"8C",x"DD",x"4E",x"FC",x"06",x"00",x"EB",x"09", -- 0x0D78
    x"E5",x"DD",x"6E",x"04",x"DD",x"66",x"05",x"C1", -- 0x0D80
    x"71",x"23",x"70",x"3E",x"20",x"DD",x"BE",x"FA", -- 0x0D88
    x"38",x"04",x"3E",x"01",x"18",x"01",x"AF",x"FD", -- 0x0D90
    x"77",x"0B",x"AF",x"FD",x"E1",x"C3",x"E4",x"82", -- 0x0D98
    x"CD",x"D0",x"82",x"FE",x"FF",x"FD",x"E5",x"DD", -- 0x0DA0
    x"6E",x"02",x"DD",x"66",x"03",x"E5",x"FD",x"E1", -- 0x0DA8
    x"DD",x"6E",x"08",x"DD",x"66",x"09",x"7E",x"FE", -- 0x0DB0
    x"20",x"20",x"0A",x"DD",x"34",x"08",x"20",x"F0", -- 0x0DB8
    x"DD",x"34",x"09",x"18",x"EB",x"7E",x"FE",x"2F", -- 0x0DC0
    x"20",x"08",x"DD",x"34",x"08",x"20",x"03",x"DD", -- 0x0DC8
    x"34",x"09",x"AF",x"FD",x"77",x"04",x"FD",x"77", -- 0x0DD0
    x"05",x"DD",x"6E",x"08",x"DD",x"66",x"09",x"3E", -- 0x0DD8
    x"20",x"BE",x"38",x"13",x"FD",x"E5",x"D1",x"CD", -- 0x0DE0
    x"87",x"8A",x"DD",x"77",x"FE",x"DD",x"6E",x"04", -- 0x0DE8
    x"DD",x"66",x"05",x"36",x"00",x"18",x"6D",x"21", -- 0x0DF0
    x"0C",x"00",x"39",x"4D",x"44",x"FD",x"E5",x"D1", -- 0x0DF8
    x"CD",x"9C",x"8C",x"DD",x"77",x"FE",x"B7",x"20", -- 0x0E00
    x"5B",x"DD",x"4E",x"04",x"DD",x"46",x"05",x"FD", -- 0x0E08
    x"E5",x"D1",x"CD",x"10",x"8C",x"DD",x"77",x"FE", -- 0x0E10
    x"B7",x"28",x"14",x"FE",x"03",x"20",x"45",x"FD", -- 0x0E18
    x"6E",x"02",x"FD",x"66",x"03",x"01",x"0B",x"00", -- 0x0E20
    x"09",x"7E",x"B7",x"20",x"37",x"18",x"1B",x"FD", -- 0x0E28
    x"6E",x"02",x"FD",x"66",x"03",x"01",x"0B",x"00", -- 0x0E30
    x"09",x"7E",x"B7",x"20",x"27",x"69",x"60",x"DD", -- 0x0E38
    x"4E",x"04",x"DD",x"46",x"05",x"09",x"CB",x"66", -- 0x0E40
    x"20",x"06",x"DD",x"36",x"FE",x"04",x"18",x"14", -- 0x0E48
    x"21",x"1A",x"00",x"09",x"23",x"56",x"21",x"1A", -- 0x0E50
    x"00",x"09",x"4E",x"B1",x"FD",x"77",x"04",x"FD", -- 0x0E58
    x"72",x"05",x"18",x"93",x"DD",x"7E",x"FE",x"FD", -- 0x0E60
    x"E1",x"C3",x"E4",x"82",x"C5",x"DD",x"E5",x"D5", -- 0x0E68
    x"DD",x"E1",x"21",x"02",x"00",x"E5",x"21",x"FE", -- 0x0E70
    x"01",x"E5",x"21",x"0A",x"00",x"39",x"4E",x"23", -- 0x0E78
    x"46",x"23",x"5E",x"23",x"56",x"D5",x"C5",x"DD", -- 0x0E80
    x"E5",x"D1",x"CD",x"4F",x"88",x"E1",x"E1",x"E1", -- 0x0E88
    x"E1",x"B7",x"28",x"05",x"3E",x"03",x"C3",x"1A", -- 0x0E90
    x"8F",x"DD",x"46",x"01",x"DD",x"5E",x"00",x"B3", -- 0x0E98
    x"6F",x"78",x"B7",x"67",x"01",x"55",x"AA",x"ED", -- 0x0EA0
    x"42",x"28",x"04",x"3E",x"02",x"18",x"6B",x"23", -- 0x0EA8
    x"23",x"E5",x"2E",x"36",x"E5",x"2E",x"0A",x"39", -- 0x0EB0
    x"4E",x"23",x"46",x"23",x"5E",x"23",x"56",x"D5", -- 0x0EB8
    x"C5",x"DD",x"E5",x"D1",x"CD",x"4F",x"88",x"E1", -- 0x0EC0
    x"E1",x"E1",x"E1",x"B7",x"20",x"12",x"DD",x"46", -- 0x0EC8
    x"01",x"DD",x"5E",x"00",x"B3",x"6F",x"78",x"B7", -- 0x0ED0
    x"67",x"01",x"46",x"41",x"ED",x"42",x"28",x"35", -- 0x0ED8
    x"AF",x"28",x"35",x"21",x"02",x"00",x"E5",x"2E", -- 0x0EE0
    x"52",x"E5",x"2E",x"0A",x"39",x"4E",x"23",x"46", -- 0x0EE8
    x"23",x"5E",x"23",x"56",x"D5",x"C5",x"DD",x"E5", -- 0x0EF0
    x"D1",x"CD",x"4F",x"88",x"E1",x"E1",x"E1",x"E1", -- 0x0EF8
    x"B7",x"20",x"15",x"DD",x"46",x"01",x"DD",x"5E", -- 0x0F00
    x"00",x"B3",x"6F",x"78",x"B7",x"67",x"01",x"46", -- 0x0F08
    x"41",x"ED",x"42",x"20",x"03",x"AF",x"18",x"02", -- 0x0F10
    x"3E",x"01",x"DD",x"E1",x"C1",x"C9",x"CD",x"D0", -- 0x0F18
    x"82",x"CA",x"FF",x"FD",x"E5",x"DD",x"6E",x"02", -- 0x0F20
    x"DD",x"66",x"03",x"E5",x"FD",x"E1",x"21",x"00", -- 0x0F28
    x"00",x"22",x"8E",x"70",x"FD",x"E5",x"E1",x"7D", -- 0x0F30
    x"B4",x"CA",x"3F",x"92",x"CD",x"00",x"87",x"CB", -- 0x0F38
    x"47",x"28",x"05",x"3E",x"02",x"C3",x"40",x"92", -- 0x0F40
    x"21",x"00",x"00",x"E5",x"E5",x"2E",x"18",x"39", -- 0x0F48
    x"EB",x"CD",x"6C",x"8E",x"E1",x"E1",x"DD",x"77", -- 0x0F50
    x"CA",x"AF",x"DD",x"77",x"D0",x"DD",x"77",x"D1", -- 0x0F58
    x"DD",x"77",x"D2",x"DD",x"77",x"D3",x"DD",x"46", -- 0x0F60
    x"CA",x"05",x"20",x"67",x"21",x"10",x"00",x"E5", -- 0x0F68
    x"21",x"BE",x"01",x"E5",x"6F",x"65",x"E5",x"E5", -- 0x0F70
    x"2E",x"1C",x"39",x"EB",x"CD",x"4F",x"88",x"E1", -- 0x0F78
    x"E1",x"E1",x"E1",x"B7",x"28",x"06",x"DD",x"36", -- 0x0F80
    x"CA",x"03",x"18",x"47",x"DD",x"7E",x"E0",x"B7", -- 0x0F88
    x"28",x"41",x"DD",x"6E",x"E4",x"48",x"61",x"C5", -- 0x0F90
    x"E5",x"DD",x"46",x"E5",x"4C",x"69",x"60",x"41", -- 0x0F98
    x"C5",x"E5",x"DD",x"6E",x"E6",x"61",x"44",x"4D", -- 0x0FA0
    x"6C",x"C5",x"E5",x"DD",x"46",x"E7",x"6C",x"CD", -- 0x0FA8
    x"52",x"92",x"CD",x"2D",x"82",x"CD",x"2D",x"82", -- 0x0FB0
    x"DD",x"75",x"D0",x"DD",x"74",x"D1",x"DD",x"71", -- 0x0FB8
    x"D2",x"DD",x"70",x"D3",x"C5",x"E5",x"21",x"18", -- 0x0FC0
    x"00",x"39",x"EB",x"CD",x"6C",x"8E",x"E1",x"E1", -- 0x0FC8
    x"DD",x"77",x"CA",x"DD",x"7E",x"CA",x"FE",x"03", -- 0x0FD0
    x"28",x"2B",x"AF",x"DD",x"B6",x"CA",x"C2",x"8F", -- 0x0FD8
    x"91",x"21",x"24",x"00",x"E5",x"2E",x"0D",x"E5", -- 0x0FE0
    x"DD",x"6E",x"D2",x"DD",x"66",x"D3",x"E5",x"DD", -- 0x0FE8
    x"6E",x"D0",x"DD",x"66",x"D1",x"E5",x"21",x"1C", -- 0x0FF0
    x"00",x"39",x"EB",x"CD",x"4F",x"88",x"E1",x"E1", -- 0x0FF8
    x"E1",x"E1",x"B7",x"28",x"05",x"3E",x"01",x"C3", -- 0x1000
    x"40",x"92",x"DD",x"66",x"E6",x"4F",x"51",x"DD", -- 0x1008
    x"5E",x"E5",x"79",x"B3",x"6F",x"DD",x"75",x"CC", -- 0x1010
    x"41",x"DD",x"74",x"CD",x"DD",x"71",x"CE",x"DD", -- 0x1018
    x"70",x"CF",x"7D",x"B4",x"20",x"2F",x"DD",x"6E", -- 0x1020
    x"F3",x"61",x"C5",x"E5",x"DD",x"66",x"F4",x"4A", -- 0x1028
    x"69",x"41",x"C5",x"E5",x"DD",x"6E",x"F5",x"61", -- 0x1030
    x"44",x"4D",x"6A",x"C5",x"E5",x"DD",x"46",x"F6", -- 0x1038
    x"CD",x"50",x"92",x"CD",x"2D",x"82",x"CD",x"2D", -- 0x1040
    x"82",x"DD",x"75",x"CC",x"DD",x"74",x"CD",x"DD", -- 0x1048
    x"71",x"CE",x"DD",x"70",x"CF",x"21",x"04",x"00", -- 0x1050
    x"39",x"DD",x"5E",x"DF",x"4A",x"42",x"51",x"CD", -- 0x1058
    x"62",x"82",x"DD",x"66",x"DE",x"0E",x"00",x"79", -- 0x1060
    x"DD",x"5E",x"DD",x"B3",x"6F",x"41",x"C5",x"E5", -- 0x1068
    x"DD",x"6E",x"D0",x"DD",x"66",x"D1",x"C1",x"09", -- 0x1070
    x"EB",x"DD",x"6E",x"D2",x"DD",x"66",x"D3",x"C1", -- 0x1078
    x"ED",x"4A",x"4D",x"44",x"EB",x"FD",x"75",x"08", -- 0x1080
    x"FD",x"74",x"09",x"FD",x"71",x"0A",x"FD",x"70", -- 0x1088
    x"0B",x"DD",x"46",x"DC",x"FD",x"70",x"02",x"DD", -- 0x1090
    x"66",x"E1",x"0E",x"00",x"51",x"DD",x"5E",x"E0", -- 0x1098
    x"79",x"B3",x"FD",x"77",x"04",x"FD",x"74",x"05", -- 0x10A0
    x"DD",x"66",x"E3",x"4A",x"79",x"DD",x"5E",x"E2", -- 0x10A8
    x"B3",x"6F",x"DD",x"75",x"D8",x"41",x"DD",x"74", -- 0x10B0
    x"D9",x"DD",x"71",x"DA",x"DD",x"70",x"DB",x"7D", -- 0x10B8
    x"B4",x"20",x"2F",x"DD",x"6E",x"EF",x"61",x"C5", -- 0x10C0
    x"E5",x"DD",x"66",x"F0",x"4A",x"69",x"41",x"C5", -- 0x10C8
    x"E5",x"DD",x"6E",x"F1",x"61",x"44",x"4D",x"6A", -- 0x10D0
    x"C5",x"E5",x"DD",x"46",x"F2",x"CD",x"50",x"92", -- 0x10D8
    x"CD",x"2D",x"82",x"CD",x"2D",x"82",x"DD",x"75", -- 0x10E0
    x"D8",x"DD",x"74",x"D9",x"DD",x"71",x"DA",x"DD", -- 0x10E8
    x"70",x"DB",x"FD",x"6E",x"02",x"4A",x"61",x"42", -- 0x10F0
    x"C5",x"E5",x"CD",x"45",x"92",x"D5",x"DD",x"46", -- 0x10F8
    x"DE",x"4C",x"79",x"DD",x"6E",x"DD",x"B5",x"5F", -- 0x1100
    x"78",x"B7",x"57",x"69",x"ED",x"52",x"D1",x"A7", -- 0x1108
    x"ED",x"52",x"41",x"C5",x"E5",x"DD",x"6E",x"D8", -- 0x1110
    x"DD",x"66",x"D9",x"C1",x"09",x"EB",x"DD",x"6E", -- 0x1118
    x"DA",x"DD",x"66",x"DB",x"C1",x"ED",x"4A",x"EB", -- 0x1120
    x"A7",x"DD",x"4E",x"CC",x"DD",x"46",x"CD",x"ED", -- 0x1128
    x"42",x"EB",x"DD",x"4E",x"CE",x"DD",x"46",x"CF", -- 0x1130
    x"ED",x"42",x"CD",x"58",x"92",x"C5",x"E5",x"21", -- 0x1138
    x"02",x"00",x"C1",x"09",x"EB",x"21",x"00",x"00", -- 0x1140
    x"C1",x"ED",x"4A",x"4D",x"44",x"EB",x"DD",x"75", -- 0x1148
    x"D4",x"DD",x"74",x"D5",x"DD",x"71",x"D6",x"DD", -- 0x1150
    x"70",x"D7",x"FD",x"75",x"06",x"FD",x"74",x"07", -- 0x1158
    x"DD",x"36",x"CA",x"02",x"A7",x"01",x"F7",x"0F", -- 0x1160
    x"ED",x"42",x"DD",x"6E",x"D6",x"DD",x"66",x"D7", -- 0x1168
    x"01",x"00",x"00",x"ED",x"42",x"38",x"18",x"DD", -- 0x1170
    x"6E",x"D4",x"DD",x"66",x"D5",x"01",x"F7",x"FF", -- 0x1178
    x"ED",x"42",x"DD",x"6E",x"D6",x"DD",x"66",x"D7", -- 0x1180
    x"01",x"00",x"00",x"ED",x"42",x"38",x"05",x"3E", -- 0x1188
    x"07",x"C3",x"40",x"92",x"DD",x"46",x"CA",x"FD", -- 0x1190
    x"70",x"00",x"AF",x"28",x"2D",x"78",x"FE",x"03", -- 0x1198
    x"20",x"28",x"DD",x"6E",x"FB",x"41",x"61",x"C5", -- 0x11A0
    x"E5",x"DD",x"46",x"FC",x"4C",x"69",x"60",x"41", -- 0x11A8
    x"C5",x"E5",x"DD",x"6E",x"FD",x"61",x"44",x"4D", -- 0x11B0
    x"6C",x"C5",x"E5",x"DD",x"46",x"FE",x"6C",x"CD", -- 0x11B8
    x"52",x"92",x"CD",x"2D",x"82",x"CD",x"2D",x"82", -- 0x11C0
    x"18",x"23",x"FD",x"6E",x"0A",x"FD",x"66",x"0B", -- 0x11C8
    x"E5",x"FD",x"6E",x"08",x"FD",x"66",x"09",x"E5", -- 0x11D0
    x"DD",x"6E",x"CC",x"DD",x"66",x"CD",x"C1",x"09", -- 0x11D8
    x"EB",x"DD",x"6E",x"CE",x"DD",x"66",x"CF",x"C1", -- 0x11E0
    x"ED",x"4A",x"4D",x"44",x"EB",x"FD",x"75",x"0C", -- 0x11E8
    x"FD",x"74",x"0D",x"FD",x"71",x"0E",x"FD",x"70", -- 0x11F0
    x"0F",x"CD",x"45",x"92",x"EB",x"01",x"00",x"00", -- 0x11F8
    x"C5",x"E5",x"FD",x"6E",x"08",x"FD",x"66",x"09", -- 0x1200
    x"C1",x"09",x"EB",x"FD",x"6E",x"0A",x"FD",x"66", -- 0x1208
    x"0B",x"C1",x"ED",x"4A",x"E5",x"D5",x"DD",x"6E", -- 0x1210
    x"CC",x"DD",x"66",x"CD",x"C1",x"09",x"EB",x"DD", -- 0x1218
    x"6E",x"CE",x"DD",x"66",x"CF",x"C1",x"ED",x"4A", -- 0x1220
    x"4D",x"44",x"EB",x"FD",x"75",x"10",x"FD",x"74", -- 0x1228
    x"11",x"FD",x"71",x"12",x"FD",x"70",x"13",x"FD", -- 0x1230
    x"36",x"01",x"00",x"FD",x"22",x"8E",x"70",x"AF", -- 0x1238
    x"FD",x"E1",x"C3",x"E4",x"82",x"FD",x"5E",x"04", -- 0x1240
    x"FD",x"56",x"05",x"06",x"04",x"C3",x"B6",x"80", -- 0x1248
    x"6A",x"65",x"4D",x"C3",x"2D",x"82",x"ED",x"4A", -- 0x1250
    x"4D",x"44",x"EB",x"C3",x"8F",x"81",x"CD",x"D0", -- 0x1258
    x"82",x"C6",x"FF",x"FD",x"E5",x"FD",x"2A",x"8E", -- 0x1260
    x"70",x"2A",x"8E",x"70",x"7D",x"B4",x"20",x"05", -- 0x1268
    x"3E",x"06",x"C3",x"FD",x"92",x"FD",x"36",x"01", -- 0x1270
    x"00",x"21",x"30",x"00",x"39",x"DD",x"75",x"EA", -- 0x1278
    x"DD",x"74",x"EB",x"DD",x"6E",x"02",x"DD",x"66", -- 0x1280
    x"03",x"E5",x"21",x"06",x"00",x"39",x"4D",x"44", -- 0x1288
    x"21",x"26",x"00",x"39",x"EB",x"CD",x"A0",x"8D", -- 0x1290
    x"E1",x"B7",x"20",x"61",x"DD",x"B6",x"C8",x"28", -- 0x1298
    x"06",x"DD",x"CB",x"D3",x"66",x"28",x"04",x"3E", -- 0x12A0
    x"03",x"18",x"52",x"DD",x"66",x"E3",x"0E",x"00", -- 0x12A8
    x"51",x"DD",x"5E",x"E2",x"79",x"B3",x"FD",x"77", -- 0x12B0
    x"1C",x"FD",x"74",x"1D",x"DD",x"6E",x"E4",x"41", -- 0x12B8
    x"61",x"C5",x"E5",x"DD",x"66",x"E5",x"4A",x"69", -- 0x12C0
    x"41",x"C5",x"E5",x"DD",x"6E",x"E6",x"61",x"44", -- 0x12C8
    x"4D",x"6A",x"C5",x"E5",x"DD",x"46",x"E7",x"CD", -- 0x12D0
    x"50",x"92",x"CD",x"2D",x"82",x"CD",x"2D",x"82", -- 0x12D8
    x"FD",x"75",x"18",x"FD",x"74",x"19",x"FD",x"71", -- 0x12E0
    x"1A",x"FD",x"70",x"1B",x"AF",x"FD",x"77",x"14", -- 0x12E8
    x"FD",x"77",x"15",x"FD",x"77",x"16",x"FD",x"77", -- 0x12F0
    x"17",x"FD",x"36",x"01",x"01",x"FD",x"E1",x"C3", -- 0x12F8
    x"E4",x"82",x"CD",x"D0",x"82",x"F0",x"FF",x"FD", -- 0x1300
    x"E5",x"DD",x"6E",x"02",x"DD",x"66",x"03",x"DD", -- 0x1308
    x"75",x"F2",x"DD",x"74",x"F3",x"FD",x"2A",x"8E", -- 0x1310
    x"70",x"DD",x"6E",x"08",x"DD",x"66",x"09",x"AF", -- 0x1318
    x"77",x"23",x"77",x"FD",x"E5",x"E1",x"7D",x"B4", -- 0x1320
    x"20",x"05",x"3E",x"06",x"C3",x"D9",x"94",x"FD", -- 0x1328
    x"CB",x"01",x"46",x"20",x"05",x"3E",x"05",x"C3", -- 0x1330
    x"D9",x"94",x"FD",x"6E",x"18",x"FD",x"66",x"19", -- 0x1338
    x"FD",x"4E",x"14",x"FD",x"46",x"15",x"ED",x"42", -- 0x1340
    x"EB",x"FD",x"6E",x"1A",x"FD",x"66",x"1B",x"FD", -- 0x1348
    x"4E",x"16",x"FD",x"46",x"17",x"ED",x"42",x"4D", -- 0x1350
    x"44",x"EB",x"DD",x"75",x"F4",x"DD",x"74",x"F5", -- 0x1358
    x"DD",x"71",x"F6",x"DD",x"70",x"F7",x"DD",x"5E", -- 0x1360
    x"04",x"DD",x"56",x"05",x"01",x"00",x"00",x"C5", -- 0x1368
    x"D5",x"A7",x"C1",x"ED",x"42",x"DD",x"6E",x"F6", -- 0x1370
    x"DD",x"66",x"F7",x"C1",x"ED",x"42",x"30",x"0C", -- 0x1378
    x"DD",x"6E",x"F4",x"DD",x"66",x"F5",x"DD",x"75", -- 0x1380
    x"04",x"DD",x"74",x"05",x"DD",x"7E",x"04",x"DD", -- 0x1388
    x"B6",x"05",x"CA",x"D9",x"94",x"FD",x"6E",x"14", -- 0x1390
    x"FD",x"7E",x"15",x"E6",x"01",x"67",x"7D",x"B4", -- 0x1398
    x"C2",x"27",x"94",x"CD",x"DE",x"94",x"FD",x"7E", -- 0x13A0
    x"02",x"C6",x"FF",x"A5",x"DD",x"77",x"FE",x"20", -- 0x13A8
    x"30",x"FD",x"7E",x"14",x"FD",x"B6",x"15",x"FD", -- 0x13B0
    x"B6",x"16",x"FD",x"B6",x"17",x"20",x"08",x"FD", -- 0x13B8
    x"6E",x"1C",x"FD",x"66",x"1D",x"18",x"09",x"FD", -- 0x13C0
    x"5E",x"1E",x"FD",x"56",x"1F",x"CD",x"B5",x"89", -- 0x13C8
    x"4D",x"44",x"21",x"01",x"00",x"A7",x"ED",x"42", -- 0x13D0
    x"D2",x"D3",x"94",x"FD",x"71",x"1E",x"FD",x"70", -- 0x13D8
    x"1F",x"FD",x"5E",x"1E",x"FD",x"56",x"1F",x"CD", -- 0x13E0
    x"2C",x"8A",x"DD",x"75",x"F8",x"DD",x"74",x"F9", -- 0x13E8
    x"DD",x"71",x"FA",x"DD",x"70",x"FB",x"7D",x"B4", -- 0x13F0
    x"B1",x"B0",x"CA",x"D3",x"94",x"DD",x"6E",x"FE", -- 0x13F8
    x"01",x"00",x"00",x"61",x"C5",x"E5",x"DD",x"6E", -- 0x1400
    x"F8",x"DD",x"66",x"F9",x"C1",x"09",x"EB",x"DD", -- 0x1408
    x"6E",x"FA",x"DD",x"66",x"FB",x"C1",x"ED",x"4A", -- 0x1410
    x"4D",x"44",x"EB",x"FD",x"75",x"20",x"FD",x"74", -- 0x1418
    x"21",x"FD",x"71",x"22",x"FD",x"70",x"23",x"FD", -- 0x1420
    x"4E",x"14",x"FD",x"7E",x"15",x"E6",x"01",x"47", -- 0x1428
    x"21",x"00",x"02",x"ED",x"42",x"DD",x"75",x"F0", -- 0x1430
    x"DD",x"74",x"F1",x"4D",x"44",x"DD",x"6E",x"04", -- 0x1438
    x"DD",x"66",x"05",x"A7",x"ED",x"42",x"30",x"0C", -- 0x1440
    x"DD",x"6E",x"04",x"DD",x"66",x"05",x"DD",x"75", -- 0x1448
    x"F0",x"DD",x"74",x"F1",x"DD",x"6E",x"F0",x"DD", -- 0x1450
    x"66",x"F1",x"E5",x"FD",x"6E",x"14",x"FD",x"7E", -- 0x1458
    x"15",x"E6",x"01",x"67",x"E5",x"FD",x"6E",x"22", -- 0x1460
    x"FD",x"66",x"23",x"E5",x"FD",x"6E",x"20",x"FD", -- 0x1468
    x"66",x"21",x"E5",x"DD",x"7E",x"02",x"DD",x"B6", -- 0x1470
    x"03",x"20",x"04",x"5F",x"57",x"18",x"06",x"DD", -- 0x1478
    x"5E",x"F2",x"DD",x"56",x"F3",x"CD",x"4F",x"88", -- 0x1480
    x"E1",x"E1",x"E1",x"E1",x"B7",x"20",x"44",x"21", -- 0x1488
    x"14",x"00",x"FD",x"E5",x"C1",x"09",x"DD",x"5E", -- 0x1490
    x"F0",x"DD",x"56",x"F1",x"4F",x"47",x"CD",x"7B", -- 0x1498
    x"82",x"21",x"04",x"00",x"39",x"7E",x"DD",x"86", -- 0x14A0
    x"F0",x"77",x"23",x"7E",x"DD",x"8E",x"F1",x"77", -- 0x14A8
    x"21",x"16",x"00",x"39",x"7E",x"DD",x"96",x"F0", -- 0x14B0
    x"77",x"23",x"7E",x"DD",x"9E",x"F1",x"77",x"DD", -- 0x14B8
    x"6E",x"08",x"DD",x"66",x"09",x"7E",x"DD",x"86", -- 0x14C0
    x"F0",x"77",x"23",x"7E",x"DD",x"8E",x"F1",x"77", -- 0x14C8
    x"C3",x"8C",x"93",x"FD",x"36",x"01",x"00",x"3E", -- 0x14D0
    x"01",x"FD",x"E1",x"C3",x"E4",x"82",x"FD",x"4E", -- 0x14D8
    x"16",x"FD",x"46",x"17",x"FD",x"6E",x"14",x"FD", -- 0x14E0
    x"66",x"15",x"3E",x"09",x"C3",x"0C",x"81",x"CD", -- 0x14E8
    x"D0",x"82",x"F2",x"FF",x"FD",x"E5",x"FD",x"2A", -- 0x14F0
    x"8E",x"70",x"2A",x"8E",x"70",x"7D",x"B4",x"20", -- 0x14F8
    x"05",x"3E",x"06",x"C3",x"5F",x"97",x"FD",x"CB", -- 0x1500
    x"01",x"46",x"20",x"05",x"3E",x"05",x"C3",x"5F", -- 0x1508
    x"97",x"FD",x"6E",x"18",x"FD",x"66",x"19",x"DD", -- 0x1510
    x"4E",x"02",x"DD",x"46",x"03",x"ED",x"42",x"FD", -- 0x1518
    x"6E",x"1A",x"FD",x"66",x"1B",x"DD",x"4E",x"04", -- 0x1520
    x"DD",x"46",x"05",x"ED",x"42",x"30",x"18",x"FD", -- 0x1528
    x"4E",x"1A",x"FD",x"46",x"1B",x"FD",x"6E",x"18", -- 0x1530
    x"DD",x"75",x"02",x"FD",x"66",x"19",x"DD",x"74", -- 0x1538
    x"03",x"DD",x"71",x"04",x"DD",x"70",x"05",x"FD", -- 0x1540
    x"4E",x"16",x"FD",x"46",x"17",x"FD",x"6E",x"14", -- 0x1548
    x"DD",x"75",x"F8",x"FD",x"66",x"15",x"DD",x"74", -- 0x1550
    x"F9",x"DD",x"71",x"FA",x"DD",x"70",x"FB",x"AF", -- 0x1558
    x"FD",x"77",x"14",x"FD",x"77",x"15",x"FD",x"77", -- 0x1560
    x"16",x"FD",x"77",x"17",x"DD",x"7E",x"02",x"DD", -- 0x1568
    x"B6",x"03",x"DD",x"B6",x"04",x"DD",x"B6",x"05", -- 0x1570
    x"CA",x"56",x"97",x"FD",x"6E",x"02",x"01",x"00", -- 0x1578
    x"00",x"61",x"3E",x"09",x"CD",x"F4",x"80",x"DD", -- 0x1580
    x"75",x"F4",x"DD",x"74",x"F5",x"DD",x"71",x"F6", -- 0x1588
    x"DD",x"70",x"F7",x"DD",x"7E",x"F8",x"DD",x"B6", -- 0x1590
    x"F9",x"DD",x"B6",x"FA",x"DD",x"B6",x"FB",x"CA", -- 0x1598
    x"59",x"96",x"C5",x"E5",x"21",x"FF",x"FF",x"E5", -- 0x15A0
    x"E5",x"DD",x"6E",x"F8",x"DD",x"66",x"F9",x"C1", -- 0x15A8
    x"09",x"EB",x"DD",x"6E",x"FA",x"DD",x"66",x"FB", -- 0x15B0
    x"C1",x"CD",x"56",x"92",x"C5",x"E5",x"DD",x"6E", -- 0x15B8
    x"F6",x"DD",x"66",x"F7",x"E5",x"DD",x"6E",x"F4", -- 0x15C0
    x"DD",x"66",x"F5",x"E5",x"21",x"FF",x"FF",x"E5", -- 0x15C8
    x"E5",x"DD",x"6E",x"02",x"DD",x"66",x"03",x"C1", -- 0x15D0
    x"09",x"EB",x"DD",x"6E",x"04",x"DD",x"66",x"05", -- 0x15D8
    x"C1",x"CD",x"56",x"92",x"59",x"50",x"A7",x"C1", -- 0x15E0
    x"ED",x"42",x"EB",x"C1",x"ED",x"42",x"38",x"69", -- 0x15E8
    x"21",x"FF",x"FF",x"E5",x"E5",x"DD",x"6E",x"F4", -- 0x15F0
    x"DD",x"66",x"F5",x"C1",x"09",x"EB",x"DD",x"6E", -- 0x15F8
    x"F6",x"DD",x"66",x"F7",x"C1",x"ED",x"4A",x"4D", -- 0x1600
    x"44",x"EB",x"CD",x"53",x"82",x"C5",x"E5",x"21", -- 0x1608
    x"FF",x"FF",x"E5",x"E5",x"DD",x"6E",x"F8",x"DD", -- 0x1610
    x"66",x"F9",x"C1",x"09",x"EB",x"DD",x"6E",x"FA", -- 0x1618
    x"DD",x"66",x"FB",x"C1",x"ED",x"4A",x"4D",x"44", -- 0x1620
    x"EB",x"CD",x"0F",x"82",x"FD",x"75",x"14",x"FD", -- 0x1628
    x"74",x"15",x"FD",x"71",x"16",x"FD",x"70",x"17", -- 0x1630
    x"21",x"12",x"00",x"39",x"FD",x"4E",x"16",x"FD", -- 0x1638
    x"46",x"17",x"FD",x"5E",x"14",x"FD",x"56",x"15", -- 0x1640
    x"CD",x"94",x"82",x"FD",x"6E",x"1E",x"DD",x"75", -- 0x1648
    x"F2",x"FD",x"66",x"1F",x"DD",x"74",x"F3",x"18", -- 0x1650
    x"12",x"FD",x"6E",x"1C",x"DD",x"75",x"F2",x"FD", -- 0x1658
    x"66",x"1D",x"DD",x"74",x"F3",x"FD",x"75",x"1E", -- 0x1660
    x"FD",x"74",x"1F",x"A7",x"DD",x"6E",x"F4",x"DD", -- 0x1668
    x"66",x"F5",x"DD",x"4E",x"02",x"DD",x"46",x"03", -- 0x1670
    x"ED",x"42",x"DD",x"6E",x"F6",x"DD",x"66",x"F7", -- 0x1678
    x"DD",x"4E",x"04",x"DD",x"46",x"05",x"ED",x"42", -- 0x1680
    x"30",x"65",x"DD",x"5E",x"F2",x"DD",x"56",x"F3", -- 0x1688
    x"CD",x"B5",x"89",x"DD",x"75",x"F2",x"DD",x"74", -- 0x1690
    x"F3",x"4D",x"44",x"21",x"01",x"00",x"A7",x"ED", -- 0x1698
    x"42",x"30",x"11",x"FD",x"4E",x"06",x"FD",x"46", -- 0x16A0
    x"07",x"DD",x"6E",x"F2",x"DD",x"66",x"F3",x"A7", -- 0x16A8
    x"ED",x"42",x"38",x"03",x"C3",x"59",x"97",x"DD", -- 0x16B0
    x"6E",x"F2",x"FD",x"75",x"1E",x"DD",x"66",x"F3", -- 0x16B8
    x"FD",x"74",x"1F",x"21",x"14",x"00",x"FD",x"E5", -- 0x16C0
    x"C1",x"09",x"DD",x"4E",x"F6",x"DD",x"46",x"F7", -- 0x16C8
    x"DD",x"5E",x"F4",x"DD",x"56",x"F5",x"CD",x"7B", -- 0x16D0
    x"82",x"21",x"12",x"00",x"39",x"DD",x"4E",x"F6", -- 0x16D8
    x"DD",x"46",x"F7",x"DD",x"5E",x"F4",x"DD",x"56", -- 0x16E0
    x"F5",x"CD",x"94",x"82",x"C3",x"6B",x"96",x"21", -- 0x16E8
    x"14",x"00",x"FD",x"E5",x"C1",x"09",x"DD",x"4E", -- 0x16F0
    x"04",x"DD",x"46",x"05",x"DD",x"5E",x"02",x"DD", -- 0x16F8
    x"56",x"03",x"CD",x"7B",x"82",x"DD",x"5E",x"F2", -- 0x1700
    x"DD",x"56",x"F3",x"CD",x"2C",x"8A",x"DD",x"75", -- 0x1708
    x"FC",x"DD",x"74",x"FD",x"DD",x"71",x"FE",x"DD", -- 0x1710
    x"70",x"FF",x"7D",x"B4",x"B1",x"B0",x"28",x"39", -- 0x1718
    x"FD",x"6E",x"02",x"26",x"00",x"2B",x"7C",x"07", -- 0x1720
    x"9F",x"4F",x"41",x"C5",x"E5",x"CD",x"DE",x"94", -- 0x1728
    x"CD",x"0F",x"82",x"C5",x"E5",x"DD",x"6E",x"FC", -- 0x1730
    x"DD",x"66",x"FD",x"C1",x"09",x"EB",x"DD",x"6E", -- 0x1738
    x"FE",x"DD",x"66",x"FF",x"C1",x"ED",x"4A",x"4D", -- 0x1740
    x"44",x"EB",x"FD",x"75",x"20",x"FD",x"74",x"21", -- 0x1748
    x"FD",x"71",x"22",x"FD",x"70",x"23",x"AF",x"18", -- 0x1750
    x"06",x"FD",x"36",x"01",x"00",x"3E",x"01",x"FD", -- 0x1758
    x"E1",x"C3",x"E4",x"82",x"CD",x"C4",x"82",x"DD", -- 0x1760
    x"56",x"04",x"DD",x"5E",x"02",x"CD",x"8B",x"97", -- 0x1768
    x"D5",x"DD",x"5E",x"08",x"DD",x"56",x"09",x"CD", -- 0x1770
    x"94",x"97",x"06",x"00",x"4D",x"DD",x"6E",x"08", -- 0x1778
    x"DD",x"66",x"09",x"D1",x"79",x"CD",x"DF",x"1F", -- 0x1780
    x"C3",x"E4",x"82",x"CD",x"C0",x"08",x"2A",x"F6", -- 0x1788
    x"73",x"19",x"EB",x"C9",x"21",x"00",x"00",x"1A", -- 0x1790
    x"B7",x"C8",x"23",x"13",x"18",x"F9",x"CD",x"C4", -- 0x1798
    x"82",x"51",x"CD",x"E8",x"85",x"DD",x"6E",x"08", -- 0x17A0
    x"DD",x"66",x"09",x"DD",x"4E",x"0A",x"DD",x"46", -- 0x17A8
    x"0B",x"CD",x"DF",x"1F",x"C3",x"E4",x"82",x"CD", -- 0x17B0
    x"C4",x"82",x"CD",x"76",x"1F",x"DD",x"66",x"02", -- 0x17B8
    x"2E",x"00",x"CD",x"79",x"1F",x"E5",x"DD",x"66", -- 0x17C0
    x"02",x"2E",x"01",x"CD",x"79",x"1F",x"7C",x"17", -- 0x17C8
    x"E1",x"B4",x"67",x"C3",x"E4",x"82",x"DD",x"E5", -- 0x17D0
    x"3A",x"C4",x"73",x"F6",x"40",x"4F",x"06",x"01", -- 0x17D8
    x"CD",x"D9",x"1F",x"DD",x"E1",x"C9",x"CD",x"C4", -- 0x17E0
    x"82",x"DD",x"7E",x"02",x"21",x"00",x"20",x"11", -- 0x17E8
    x"20",x"00",x"CD",x"82",x"1F",x"C3",x"E4",x"82", -- 0x17F0
    x"DD",x"E5",x"CD",x"85",x"1F",x"DD",x"E1",x"C9", -- 0x17F8
    x"DD",x"E5",x"CD",x"E9",x"18",x"DD",x"E1",x"C9", -- 0x1800
    x"3D",x"3E",x"00",x"45",x"72",x"72",x"6F",x"72", -- 0x1808
    x"2E",x"2E",x"2E",x"2E",x"2E",x"2E",x"52",x"65", -- 0x1810
    x"73",x"65",x"74",x"00",x"4D",x"45",x"4E",x"55", -- 0x1818
    x"2E",x"54",x"58",x"54",x"00",x"4C",x"2D",x"46", -- 0x1820
    x"69",x"72",x"65",x"3A",x"4C",x"6F",x"61",x"64", -- 0x1828
    x"20",x"20",x"52",x"2D",x"46",x"69",x"72",x"65", -- 0x1830
    x"3A",x"52",x"65",x"73",x"74",x"61",x"72",x"74", -- 0x1838
    x"00",x"20",x"20",x"20",x"55",x"2F",x"44",x"3A", -- 0x1840
    x"53",x"65",x"6C",x"65",x"63",x"74",x"20",x"20", -- 0x1848
    x"20",x"4C",x"2F",x"52",x"3A",x"50",x"61",x"67", -- 0x1850
    x"65",x"00",x"3C",x"45",x"53",x"43",x"3E",x"52", -- 0x1858
    x"65",x"73",x"65",x"74",x"20",x"3C",x"55",x"2F", -- 0x1860
    x"44",x"3E",x"53",x"65",x"6C",x"20",x"3C",x"4C", -- 0x1868
    x"2F",x"52",x"3E",x"50",x"61",x"67",x"65",x"00", -- 0x1870
    x"3C",x"51",x"3E",x"2A",x"20",x"3C",x"57",x"3E", -- 0x1878
    x"23",x"20",x"3C",x"5A",x"3E",x"4C",x"2D",x"46", -- 0x1880
    x"69",x"72",x"65",x"20",x"3C",x"58",x"3E",x"52", -- 0x1888
    x"2D",x"46",x"69",x"72",x"65",x"00",x"20",x"20", -- 0x1890
    x"00",x"2E",x"72",x"6F",x"6D",x"00",x"4C",x"6F", -- 0x1898
    x"61",x"64",x"69",x"6E",x"67",x"00",x"43",x"6F", -- 0x18A0
    x"6C",x"65",x"63",x"6F",x"2F",x"00",x"00",x"00", -- 0x18A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1900
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1908
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1910
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1918
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1920
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1928
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1930
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1938
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1940
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1948
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1950
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1958
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1960
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1968
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1970
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1978
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1980
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1988
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1990
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1998
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x1FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
