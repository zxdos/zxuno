-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity cart_rom4 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of cart_rom4 is


  type ROM_ARRAY is array(6144 to 8191) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"A0",x"90",x"00",x"00",x"00",x"80",x"80",x"80", -- 0x0000
    x"80",x"F8",x"00",x"00",x"00",x"88",x"D8",x"A8", -- 0x0008
    x"88",x"88",x"00",x"00",x"00",x"88",x"C8",x"A8", -- 0x0010
    x"98",x"88",x"00",x"00",x"00",x"F8",x"88",x"88", -- 0x0018
    x"88",x"F8",x"00",x"00",x"00",x"F0",x"88",x"F0", -- 0x0020
    x"80",x"80",x"00",x"00",x"00",x"F8",x"88",x"A8", -- 0x0028
    x"90",x"E0",x"00",x"00",x"00",x"F8",x"88",x"F8", -- 0x0030
    x"A0",x"90",x"00",x"00",x"00",x"78",x"80",x"70", -- 0x0038
    x"08",x"F0",x"00",x"00",x"00",x"F8",x"20",x"20", -- 0x0040
    x"20",x"20",x"00",x"00",x"00",x"88",x"88",x"88", -- 0x0048
    x"88",x"70",x"00",x"00",x"00",x"88",x"88",x"90", -- 0x0050
    x"A0",x"40",x"00",x"00",x"00",x"88",x"88",x"A8", -- 0x0058
    x"D8",x"88",x"00",x"00",x"00",x"88",x"50",x"20", -- 0x0060
    x"50",x"88",x"00",x"00",x"00",x"88",x"50",x"20", -- 0x0068
    x"20",x"20",x"00",x"00",x"00",x"F8",x"10",x"20", -- 0x0070
    x"40",x"F8",x"00",x"38",x"40",x"20",x"C0",x"20", -- 0x0078
    x"40",x"38",x"00",x"40",x"20",x"10",x"08",x"10", -- 0x0080
    x"20",x"40",x"00",x"E0",x"10",x"20",x"18",x"20", -- 0x0088
    x"10",x"E0",x"00",x"40",x"A8",x"10",x"00",x"00", -- 0x0090
    x"00",x"00",x"00",x"A8",x"50",x"A8",x"50",x"A8", -- 0x0098
    x"50",x"A8",x"00",x"01",x"02",x"0E",x"0F",x"08", -- 0x00A0
    x"09",x"12",x"13",x"03",x"04",x"0E",x"0F",x"05", -- 0x00A8
    x"14",x"00",x"00",x"05",x"00",x"10",x"11",x"0A", -- 0x00B0
    x"0B",x"15",x"16",x"06",x"07",x"10",x"11",x"05", -- 0x00B8
    x"14",x"00",x"00",x"01",x"02",x"0E",x"0F",x"03", -- 0x00C0
    x"04",x"0E",x"0F",x"03",x"04",x"0E",x"0F",x"0C", -- 0x00C8
    x"0D",x"17",x"18",x"FF",x"4F",x"7D",x"D3",x"BF", -- 0x00D0
    x"7C",x"F6",x"40",x"D3",x"BF",x"79",x"D3",x"BE", -- 0x00D8
    x"1B",x"7A",x"B3",x"20",x"F8",x"CD",x"DC",x"1F", -- 0x00E0
    x"C9",x"06",x"00",x"0E",x"00",x"CD",x"D9",x"1F", -- 0x00E8
    x"06",x"01",x"0E",x"80",x"CD",x"D9",x"1F",x"3E", -- 0x00F0
    x"02",x"21",x"00",x"18",x"CD",x"B8",x"1F",x"3E", -- 0x00F8
    x"04",x"21",x"00",x"20",x"CD",x"B8",x"1F",x"3E", -- 0x0100
    x"03",x"21",x"00",x"00",x"CD",x"B8",x"1F",x"3E", -- 0x0108
    x"00",x"21",x"00",x"1B",x"CD",x"B8",x"1F",x"3E", -- 0x0110
    x"01",x"21",x"00",x"38",x"CD",x"B8",x"1F",x"06", -- 0x0118
    x"07",x"0E",x"00",x"CD",x"D9",x"1F",x"C9",x"21", -- 0x0120
    x"8B",x"15",x"11",x"1D",x"00",x"FD",x"21",x"60", -- 0x0128
    x"00",x"3E",x"03",x"CD",x"BE",x"1F",x"21",x"A3", -- 0x0130
    x"15",x"11",x"00",x"00",x"FD",x"21",x"01",x"00", -- 0x0138
    x"3E",x"03",x"CD",x"BE",x"1F",x"C9",x"01",x"00", -- 0x0140
    x"00",x"7E",x"FE",x"2F",x"C8",x"23",x"03",x"18", -- 0x0148
    x"F8",x"C5",x"FD",x"E1",x"3E",x"20",x"99",x"1F", -- 0x0150
    x"06",x"00",x"4F",x"09",x"44",x"4D",x"62",x"6B", -- 0x0158
    x"50",x"59",x"3E",x"02",x"CD",x"BE",x"1F",x"C9", -- 0x0160
    x"21",x"00",x"17",x"11",x"FF",x"00",x"1B",x"7A", -- 0x0168
    x"B3",x"20",x"FB",x"2B",x"7C",x"B5",x"20",x"F3", -- 0x0170
    x"C9",x"21",x"00",x"00",x"11",x"00",x"40",x"3E", -- 0x0178
    x"00",x"CD",x"82",x"1F",x"CD",x"85",x"1F",x"06", -- 0x0180
    x"0F",x"0E",x"04",x"CD",x"D9",x"1F",x"CD",x"7F", -- 0x0188
    x"1F",x"21",x"7C",x"1A",x"11",x"25",x"00",x"FD", -- 0x0190
    x"21",x"16",x"00",x"3E",x"02",x"CD",x"BE",x"1F", -- 0x0198
    x"21",x"92",x"1A",x"11",x"65",x"00",x"FD",x"21", -- 0x01A0
    x"17",x"00",x"3E",x"02",x"CD",x"BE",x"1F",x"11", -- 0x01A8
    x"C5",x"00",x"CD",x"CA",x"1A",x"11",x"05",x"01", -- 0x01B0
    x"CD",x"CA",x"1A",x"11",x"45",x"01",x"CD",x"CA", -- 0x01B8
    x"1A",x"11",x"85",x"01",x"CD",x"CA",x"1A",x"11", -- 0x01C0
    x"E5",x"01",x"CD",x"CA",x"1A",x"11",x"25",x"02", -- 0x01C8
    x"CD",x"CA",x"1A",x"11",x"65",x"02",x"CD",x"CA", -- 0x01D0
    x"1A",x"11",x"A5",x"02",x"CD",x"CA",x"1A",x"11", -- 0x01D8
    x"05",x"01",x"CD",x"D7",x"1A",x"11",x"45",x"01", -- 0x01E0
    x"CD",x"DC",x"1A",x"11",x"85",x"01",x"CD",x"E1", -- 0x01E8
    x"1A",x"21",x"C2",x"1A",x"11",x"E5",x"01",x"CD", -- 0x01F0
    x"E4",x"1A",x"21",x"C3",x"1A",x"11",x"25",x"02", -- 0x01F8
    x"CD",x"E4",x"1A",x"21",x"C4",x"1A",x"11",x"65", -- 0x0200
    x"02",x"CD",x"E4",x"1A",x"21",x"C5",x"1A",x"11", -- 0x0208
    x"A5",x"02",x"CD",x"E4",x"1A",x"11",x"0F",x"01", -- 0x0210
    x"CD",x"D7",x"1A",x"11",x"4F",x"01",x"CD",x"DC", -- 0x0218
    x"1A",x"11",x"8F",x"01",x"CD",x"E1",x"1A",x"11", -- 0x0220
    x"F1",x"01",x"CD",x"EE",x"1A",x"11",x"31",x"02", -- 0x0228
    x"CD",x"EE",x"1A",x"11",x"71",x"02",x"CD",x"EE", -- 0x0230
    x"1A",x"11",x"B1",x"02",x"CD",x"EE",x"1A",x"11", -- 0x0238
    x"2F",x"02",x"CD",x"D7",x"1A",x"11",x"6F",x"02", -- 0x0240
    x"CD",x"DC",x"1A",x"11",x"AF",x"02",x"CD",x"E1", -- 0x0248
    x"1A",x"11",x"FB",x"01",x"CD",x"FB",x"1A",x"11", -- 0x0250
    x"3B",x"02",x"CD",x"FB",x"1A",x"11",x"7B",x"02", -- 0x0258
    x"CD",x"FB",x"1A",x"11",x"BB",x"02",x"CD",x"FB", -- 0x0260
    x"1A",x"2A",x"FA",x"73",x"11",x"20",x"00",x"3E", -- 0x0268
    x"F4",x"CD",x"82",x"1F",x"06",x"01",x"0E",x"C0", -- 0x0270
    x"CD",x"D9",x"1F",x"C9",x"54",x"4F",x"20",x"53", -- 0x0278
    x"45",x"4C",x"45",x"43",x"54",x"20",x"47",x"41", -- 0x0280
    x"4D",x"45",x"20",x"4F",x"50",x"54",x"49",x"4F", -- 0x0288
    x"4E",x"2C",x"50",x"52",x"45",x"53",x"53",x"20", -- 0x0290
    x"42",x"55",x"54",x"54",x"4F",x"4E",x"20",x"4F", -- 0x0298
    x"4E",x"20",x"4B",x"45",x"59",x"50",x"41",x"44", -- 0x02A0
    x"2E",x"31",x"20",x"3D",x"20",x"53",x"4B",x"49", -- 0x02A8
    x"4C",x"4C",x"20",x"31",x"2F",x"4F",x"4E",x"45", -- 0x02B0
    x"20",x"50",x"4C",x"41",x"59",x"45",x"52",x"32", -- 0x02B8
    x"33",x"34",x"35",x"36",x"37",x"38",x"54",x"57", -- 0x02C0
    x"4F",x"53",x"21",x"A9",x"1A",x"FD",x"21",x"16", -- 0x02C8
    x"00",x"3E",x"02",x"CD",x"BE",x"1F",x"C9",x"21", -- 0x02D0
    x"BF",x"1A",x"18",x"08",x"21",x"C0",x"1A",x"18", -- 0x02D8
    x"03",x"21",x"C1",x"1A",x"FD",x"21",x"01",x"00", -- 0x02E0
    x"3E",x"02",x"CD",x"BE",x"1F",x"C9",x"21",x"C6", -- 0x02E8
    x"1A",x"FD",x"21",x"03",x"00",x"3E",x"02",x"CD", -- 0x02F0
    x"BE",x"1F",x"C9",x"21",x"C9",x"1A",x"FD",x"21", -- 0x02F8
    x"01",x"00",x"3E",x"02",x"CD",x"BE",x"1F",x"C9", -- 0x0300
    x"02",x"00",x"01",x"00",x"02",x"00",x"01",x"08", -- 0x0308
    x"1B",x"11",x"BA",x"73",x"CD",x"98",x"00",x"3A", -- 0x0310
    x"BA",x"73",x"2A",x"BB",x"73",x"4F",x"06",x"00", -- 0x0318
    x"DD",x"21",x"F2",x"73",x"DD",x"09",x"DD",x"09", -- 0x0320
    x"DD",x"75",x"00",x"DD",x"74",x"01",x"3A",x"C3", -- 0x0328
    x"73",x"CB",x"4F",x"28",x"27",x"79",x"FE",x"03", -- 0x0330
    x"28",x"06",x"FE",x"04",x"28",x"10",x"18",x"1C", -- 0x0338
    x"06",x"04",x"7D",x"B4",x"20",x"04",x"0E",x"03", -- 0x0340
    x"18",x"28",x"0E",x"07",x"18",x"24",x"06",x"03", -- 0x0348
    x"7D",x"B4",x"20",x"04",x"0E",x"7F",x"18",x"1A", -- 0x0350
    x"0E",x"FF",x"18",x"16",x"FD",x"21",x"76",x"1B", -- 0x0358
    x"FD",x"09",x"FD",x"09",x"FD",x"7E",x"00",x"FD", -- 0x0360
    x"46",x"01",x"CB",x"3C",x"CB",x"1D",x"3D",x"20", -- 0x0368
    x"F9",x"4D",x"CD",x"CA",x"1C",x"C9",x"07",x"05", -- 0x0370
    x"0B",x"06",x"0A",x"02",x"0B",x"04",x"06",x"03", -- 0x0378
    x"05",x"00",x"01",x"00",x"01",x"00",x"01",x"00", -- 0x0380
    x"FE",x"FF",x"02",x"00",x"01",x"80",x"1B",x"11", -- 0x0388
    x"BA",x"73",x"CD",x"98",x"00",x"3A",x"BA",x"73", -- 0x0390
    x"ED",x"5B",x"BB",x"73",x"FD",x"2A",x"BF",x"73", -- 0x0398
    x"2A",x"BD",x"73",x"CD",x"AA",x"1B",x"CD",x"3E", -- 0x03A0
    x"1D",x"C9",x"FD",x"22",x"FE",x"73",x"DD",x"21", -- 0x03A8
    x"F2",x"73",x"4F",x"06",x"00",x"FE",x"04",x"20", -- 0x03B0
    x"07",x"3A",x"C3",x"73",x"CB",x"4F",x"28",x"2C", -- 0x03B8
    x"FD",x"21",x"FF",x"1B",x"FD",x"09",x"FD",x"7E", -- 0x03C0
    x"00",x"FE",x"00",x"28",x"1F",x"CB",x"23",x"CB", -- 0x03C8
    x"12",x"3D",x"20",x"F9",x"C5",x"ED",x"4B",x"FE", -- 0x03D0
    x"73",x"FD",x"7E",x"00",x"FE",x"00",x"28",x"0B", -- 0x03D8
    x"CB",x"21",x"CB",x"10",x"3D",x"20",x"F9",x"ED", -- 0x03E0
    x"43",x"FE",x"73",x"C1",x"E5",x"DD",x"09",x"DD", -- 0x03E8
    x"09",x"DD",x"6E",x"00",x"DD",x"66",x"01",x"19", -- 0x03F0
    x"EB",x"E1",x"ED",x"4B",x"FE",x"73",x"C9",x"02", -- 0x03F8
    x"03",x"00",x"03",x"03",x"05",x"00",x"01",x"00", -- 0x0400
    x"01",x"00",x"01",x"00",x"FE",x"FF",x"02",x"00", -- 0x0408
    x"01",x"04",x"1C",x"11",x"BA",x"73",x"CD",x"98", -- 0x0410
    x"00",x"3A",x"BA",x"73",x"ED",x"5B",x"BB",x"73", -- 0x0418
    x"FD",x"2A",x"BF",x"73",x"2A",x"BD",x"73",x"F5", -- 0x0420
    x"FE",x"00",x"20",x"22",x"3A",x"C7",x"73",x"FE", -- 0x0428
    x"01",x"20",x"1B",x"F1",x"E5",x"2A",x"02",x"80", -- 0x0430
    x"7B",x"CB",x"27",x"CB",x"27",x"5F",x"19",x"EB", -- 0x0438
    x"FD",x"E5",x"C1",x"79",x"CB",x"27",x"CB",x"27", -- 0x0440
    x"4F",x"E1",x"ED",x"B0",x"18",x"07",x"F1",x"CD", -- 0x0448
    x"AA",x"1B",x"CD",x"01",x"1D",x"C9",x"01",x"00", -- 0x0450
    x"01",x"00",x"01",x"56",x"1C",x"11",x"BA",x"73", -- 0x0458
    x"CD",x"98",x"00",x"3A",x"BA",x"73",x"47",x"AF", -- 0x0460
    x"2A",x"04",x"80",x"77",x"23",x"3C",x"B8",x"20", -- 0x0468
    x"FA",x"C9",x"01",x"00",x"01",x"00",x"01",x"72", -- 0x0470
    x"1C",x"11",x"BA",x"73",x"CD",x"98",x"00",x"3A", -- 0x0478
    x"BA",x"73",x"DD",x"2A",x"04",x"80",x"F5",x"FD", -- 0x0480
    x"21",x"F2",x"73",x"FD",x"5E",x"00",x"FD",x"56", -- 0x0488
    x"01",x"7B",x"D3",x"BF",x"7A",x"F6",x"40",x"D3", -- 0x0490
    x"BF",x"F1",x"2A",x"02",x"80",x"DD",x"4E",x"00", -- 0x0498
    x"DD",x"23",x"06",x"00",x"09",x"09",x"09",x"09", -- 0x04A0
    x"06",x"04",x"0E",x"BE",x"ED",x"A3",x"00",x"00", -- 0x04A8
    x"20",x"FA",x"3D",x"20",x"E5",x"C9",x"02",x"00", -- 0x04B0
    x"01",x"00",x"01",x"00",x"01",x"B6",x"1C",x"11", -- 0x04B8
    x"BA",x"73",x"CD",x"98",x"00",x"2A",x"BA",x"73", -- 0x04C0
    x"4C",x"45",x"79",x"D3",x"BF",x"78",x"C6",x"80", -- 0x04C8
    x"D3",x"BF",x"78",x"FE",x"00",x"20",x"04",x"79", -- 0x04D0
    x"32",x"C3",x"73",x"78",x"FE",x"01",x"20",x"04", -- 0x04D8
    x"79",x"32",x"C4",x"73",x"C9",x"03",x"00",x"FE", -- 0x04E0
    x"FF",x"02",x"00",x"02",x"00",x"01",x"E5",x"1C", -- 0x04E8
    x"11",x"BA",x"73",x"CD",x"98",x"00",x"2A",x"BA", -- 0x04F0
    x"73",x"ED",x"5B",x"BC",x"73",x"ED",x"4B",x"BE", -- 0x04F8
    x"73",x"E5",x"D5",x"E1",x"11",x"00",x"40",x"19", -- 0x0500
    x"7D",x"D3",x"BF",x"7C",x"D3",x"BF",x"C5",x"D1", -- 0x0508
    x"E1",x"0E",x"BE",x"43",x"ED",x"A3",x"00",x"00", -- 0x0510
    x"C2",x"14",x"1D",x"15",x"FA",x"21",x"1D",x"20", -- 0x0518
    x"F3",x"C9",x"03",x"00",x"FE",x"FF",x"02",x"00", -- 0x0520
    x"02",x"00",x"01",x"22",x"1D",x"11",x"BA",x"73", -- 0x0528
    x"CD",x"98",x"00",x"2A",x"BA",x"73",x"ED",x"5B", -- 0x0530
    x"BC",x"73",x"ED",x"4B",x"BE",x"73",x"7B",x"D3", -- 0x0538
    x"BF",x"7A",x"D3",x"BF",x"C5",x"D1",x"0E",x"BE", -- 0x0540
    x"43",x"ED",x"A2",x"00",x"00",x"C2",x"49",x"1D", -- 0x0548
    x"15",x"FA",x"56",x"1D",x"20",x"F3",x"C9",x"DB", -- 0x0550
    x"BF",x"C9",x"DD",x"21",x"96",x"1D",x"18",x"10", -- 0x0558
    x"DD",x"21",x"B7",x"1D",x"18",x"0A",x"DD",x"21", -- 0x0560
    x"E5",x"1D",x"18",x"04",x"DD",x"21",x"07",x"1E", -- 0x0568
    x"D9",x"08",x"DD",x"E5",x"08",x"F5",x"08",x"F1", -- 0x0570
    x"D9",x"D5",x"D9",x"D1",x"FD",x"21",x"01",x"00", -- 0x0578
    x"2A",x"06",x"80",x"CD",x"A3",x"1B",x"DD",x"E1", -- 0x0580
    x"DD",x"E5",x"DD",x"E9",x"13",x"0B",x"78",x"B1", -- 0x0588
    x"D9",x"20",x"E1",x"DD",x"E1",x"C9",x"2A",x"06", -- 0x0590
    x"80",x"01",x"08",x"00",x"E5",x"D1",x"09",x"EB", -- 0x0598
    x"CD",x"00",x"1F",x"CD",x"72",x"1E",x"CD",x"5D", -- 0x05A0
    x"1E",x"FE",x"01",x"20",x"06",x"CD",x"89",x"1E", -- 0x05A8
    x"CD",x"9A",x"1E",x"D9",x"23",x"18",x"D5",x"2A", -- 0x05B0
    x"06",x"80",x"01",x"08",x"00",x"E5",x"D1",x"09", -- 0x05B8
    x"EB",x"CD",x"4E",x"1F",x"CD",x"72",x"1E",x"CD", -- 0x05C0
    x"5D",x"1E",x"FE",x"01",x"20",x"13",x"CD",x"89", -- 0x05C8
    x"1E",x"2A",x"06",x"80",x"01",x"08",x"00",x"E5", -- 0x05D0
    x"D1",x"09",x"EB",x"CD",x"4E",x"1F",x"CD",x"9A", -- 0x05D8
    x"1E",x"D9",x"23",x"18",x"A7",x"2A",x"06",x"80", -- 0x05E0
    x"01",x"08",x"00",x"E5",x"D1",x"09",x"EB",x"CD", -- 0x05E8
    x"12",x"1F",x"CD",x"72",x"1E",x"CD",x"5D",x"1E", -- 0x05F0
    x"FE",x"01",x"20",x"06",x"CD",x"89",x"1E",x"CD", -- 0x05F8
    x"9A",x"1E",x"D9",x"23",x"C3",x"8C",x"1D",x"2A", -- 0x0600
    x"06",x"80",x"01",x"08",x"00",x"E5",x"D1",x"09", -- 0x0608
    x"EB",x"CD",x"AB",x"1E",x"08",x"F5",x"08",x"F1", -- 0x0610
    x"D9",x"E5",x"D9",x"D1",x"2A",x"06",x"80",x"01", -- 0x0618
    x"08",x"00",x"09",x"FD",x"21",x"04",x"00",x"CD", -- 0x0620
    x"27",x"1C",x"CD",x"5D",x"1E",x"FE",x"01",x"20", -- 0x0628
    x"24",x"CD",x"89",x"1E",x"2A",x"06",x"80",x"01", -- 0x0630
    x"08",x"00",x"E5",x"D1",x"09",x"EB",x"CD",x"EA", -- 0x0638
    x"1E",x"3E",x"04",x"D9",x"E5",x"D9",x"D1",x"2A", -- 0x0640
    x"06",x"80",x"01",x"08",x"00",x"09",x"FD",x"21", -- 0x0648
    x"04",x"00",x"CD",x"27",x"1C",x"D9",x"23",x"23", -- 0x0650
    x"23",x"23",x"C3",x"8C",x"1D",x"08",x"F5",x"08", -- 0x0658
    x"F1",x"FE",x"03",x"20",x"0A",x"21",x"C3",x"73", -- 0x0660
    x"CB",x"4E",x"28",x"03",x"3E",x"01",x"C9",x"3E", -- 0x0668
    x"00",x"C9",x"08",x"F5",x"08",x"F1",x"D9",x"E5", -- 0x0670
    x"D9",x"D1",x"2A",x"06",x"80",x"01",x"08",x"00", -- 0x0678
    x"09",x"FD",x"21",x"01",x"00",x"CD",x"27",x"1C", -- 0x0680
    x"C9",x"3E",x"04",x"D9",x"D5",x"D9",x"D1",x"2A", -- 0x0688
    x"06",x"80",x"FD",x"21",x"01",x"00",x"CD",x"A3", -- 0x0690
    x"1B",x"C9",x"3E",x"04",x"D9",x"E5",x"D9",x"D1", -- 0x0698
    x"2A",x"06",x"80",x"FD",x"21",x"01",x"00",x"CD", -- 0x06A0
    x"27",x"1C",x"C9",x"E5",x"DD",x"E1",x"D5",x"FD", -- 0x06A8
    x"E1",x"01",x"08",x"00",x"DD",x"7E",x"00",x"DD", -- 0x06B0
    x"23",x"57",x"1E",x"04",x"CB",x"17",x"CB",x"14", -- 0x06B8
    x"CB",x"12",x"CB",x"14",x"1D",x"20",x"F5",x"1E", -- 0x06C0
    x"04",x"CB",x"17",x"CB",x"15",x"CB",x"12",x"CB", -- 0x06C8
    x"15",x"1D",x"20",x"F5",x"FD",x"74",x"00",x"FD", -- 0x06D0
    x"75",x"10",x"FD",x"23",x"FD",x"74",x"00",x"FD", -- 0x06D8
    x"75",x"10",x"FD",x"23",x"0B",x"79",x"B0",x"20", -- 0x06E0
    x"CB",x"C9",x"01",x"10",x"00",x"E5",x"7E",x"23", -- 0x06E8
    x"12",x"13",x"12",x"13",x"0B",x"79",x"FE",x"08", -- 0x06F0
    x"20",x"01",x"E1",x"79",x"B0",x"20",x"EF",x"C9", -- 0x06F8
    x"01",x"08",x"00",x"46",x"3E",x"80",x"CB",x"10", -- 0x0700
    x"1F",x"30",x"FB",x"12",x"23",x"13",x"0D",x"20", -- 0x0708
    x"F2",x"C9",x"E5",x"DD",x"E1",x"EB",x"01",x"08", -- 0x0710
    x"00",x"DD",x"CB",x"00",x"16",x"CB",x"1E",x"DD", -- 0x0718
    x"CB",x"01",x"16",x"CB",x"1E",x"DD",x"CB",x"02", -- 0x0720
    x"16",x"CB",x"1E",x"DD",x"CB",x"03",x"16",x"CB", -- 0x0728
    x"1E",x"DD",x"CB",x"04",x"16",x"CB",x"1E",x"DD", -- 0x0730
    x"CB",x"05",x"16",x"CB",x"1E",x"DD",x"CB",x"06", -- 0x0738
    x"16",x"CB",x"1E",x"DD",x"CB",x"07",x"16",x"CB", -- 0x0740
    x"1E",x"23",x"0D",x"20",x"CC",x"C9",x"01",x"07", -- 0x0748
    x"00",x"09",x"03",x"7E",x"12",x"13",x"2B",x"0B", -- 0x0750
    x"78",x"B1",x"20",x"F7",x"C9",x"FF",x"FF",x"FF", -- 0x0758
    x"FF",x"C3",x"00",x"03",x"C3",x"88",x"04",x"C3", -- 0x0760
    x"C7",x"06",x"C3",x"5A",x"1D",x"C3",x"60",x"1D", -- 0x0768
    x"C3",x"66",x"1D",x"C3",x"6C",x"1D",x"C3",x"4A", -- 0x0770
    x"11",x"C3",x"8B",x"11",x"C3",x"79",x"19",x"C3", -- 0x0778
    x"27",x"19",x"C3",x"D4",x"18",x"C3",x"E9",x"18", -- 0x0780
    x"C3",x"6A",x"11",x"C3",x"0E",x"1B",x"C3",x"8C", -- 0x0788
    x"1B",x"C3",x"10",x"1C",x"C3",x"5A",x"1C",x"C3", -- 0x0790
    x"76",x"1C",x"C3",x"9A",x"0F",x"C3",x"B8",x"0F", -- 0x0798
    x"C3",x"44",x"10",x"C3",x"BF",x"10",x"C3",x"BC", -- 0x07A0
    x"1C",x"C3",x"ED",x"1C",x"C3",x"2A",x"1D",x"C3", -- 0x07A8
    x"55",x"06",x"C3",x"03",x"02",x"C3",x"51",x"02", -- 0x07B0
    x"C3",x"1D",x"1B",x"C3",x"A3",x"1B",x"C3",x"27", -- 0x07B8
    x"1C",x"C3",x"66",x"1C",x"C3",x"82",x"1C",x"C3", -- 0x07C0
    x"AA",x"0F",x"C3",x"C4",x"0F",x"C3",x"53",x"10", -- 0x07C8
    x"C3",x"CB",x"10",x"C3",x"37",x"0F",x"C3",x"3B", -- 0x07D0
    x"02",x"C3",x"CA",x"1C",x"C3",x"57",x"1D",x"C3", -- 0x07D8
    x"01",x"1D",x"C3",x"3E",x"1D",x"C3",x"64",x"06", -- 0x07E0
    x"C3",x"79",x"06",x"C3",x"C1",x"11",x"C3",x"13", -- 0x07E8
    x"02",x"C3",x"5E",x"02",x"C3",x"7F",x"02",x"C3", -- 0x07F0
    x"A3",x"04",x"C3",x"D8",x"06",x"C3",x"3B",x"00"  -- 0x07F8
  );

signal AR	: std_logic_vector(12 downto 0);


begin

  AR(12 downto 11) <= "11";
  process(CLK)
  begin
    if CLK'event and CLK = '1' then
      AR(10 downto 0) <= ADDR(10 downto 0);   
    end if;
  end process;

    process (AR)
	 begin
	   DATA <= ROM(to_integer(unsigned(AR)));
    end process; 

end RTL;
