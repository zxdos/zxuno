library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library UNISIM;
use UNISIM.Vcomponents.all;

entity RomSmelk3006 is
    port (
        clk  : in  std_logic;
        addr : in  std_logic_vector(13 downto 0);
        data : out std_logic_vector(7 downto 0)
        );
end;

architecture RTL of RomSmelk3006 is

    signal rom_addr : std_logic_vector(13 downto 0);

begin

    p_addr : process(addr)
    begin
        rom_addr              <= (others => '0');
        rom_addr(13 downto 0) <= addr;
    end process;

    p_rom : process
    begin
        wait until rising_edge(clk);
        data <= (others => '0');
        case rom_addr is
            when "00" & x"000" => data <= x"00";
            when "00" & x"001" => data <= x"00";
            when "00" & x"002" => data <= x"00";
            when "00" & x"003" => data <= x"4c";
            when "00" & x"004" => data <= x"55";
            when "00" & x"005" => data <= x"94";
            when "00" & x"006" => data <= x"82";
            when "00" & x"007" => data <= x"11";
            when "00" & x"008" => data <= x"5a";
            when "00" & x"009" => data <= x"53";
            when "00" & x"00a" => data <= x"50";
            when "00" & x"00b" => data <= x"49";
            when "00" & x"00c" => data <= x"00";
            when "00" & x"00d" => data <= x"30";
            when "00" & x"00e" => data <= x"2e";
            when "00" & x"00f" => data <= x"39";
            when "00" & x"010" => data <= x"30";
            when "00" & x"011" => data <= x"00";
            when "00" & x"012" => data <= x"28";
            when "00" & x"013" => data <= x"43";
            when "00" & x"014" => data <= x"29";
            when "00" & x"015" => data <= x"6c";
            when "00" & x"016" => data <= x"1e";
            when "00" & x"017" => data <= x"02";
            when "00" & x"018" => data <= x"20";
            when "00" & x"019" => data <= x"5b";
            when "00" & x"01a" => data <= x"80";
            when "00" & x"01b" => data <= x"44";
            when "00" & x"01c" => data <= x"69";
            when "00" & x"01d" => data <= x"73";
            when "00" & x"01e" => data <= x"6b";
            when "00" & x"01f" => data <= x"20";
            when "00" & x"020" => data <= x"90";
            when "00" & x"021" => data <= x"11";
            when "00" & x"022" => data <= x"20";
            when "00" & x"023" => data <= x"5b";
            when "00" & x"024" => data <= x"80";
            when "00" & x"025" => data <= x"42";
            when "00" & x"026" => data <= x"61";
            when "00" & x"027" => data <= x"64";
            when "00" & x"028" => data <= x"20";
            when "00" & x"029" => data <= x"90";
            when "00" & x"02a" => data <= x"08";
            when "00" & x"02b" => data <= x"20";
            when "00" & x"02c" => data <= x"5b";
            when "00" & x"02d" => data <= x"80";
            when "00" & x"02e" => data <= x"46";
            when "00" & x"02f" => data <= x"69";
            when "00" & x"030" => data <= x"6c";
            when "00" & x"031" => data <= x"65";
            when "00" & x"032" => data <= x"20";
            when "00" & x"033" => data <= x"85";
            when "00" & x"034" => data <= x"b3";
            when "00" & x"035" => data <= x"68";
            when "00" & x"036" => data <= x"85";
            when "00" & x"037" => data <= x"ae";
            when "00" & x"038" => data <= x"68";
            when "00" & x"039" => data <= x"85";
            when "00" & x"03a" => data <= x"af";
            when "00" & x"03b" => data <= x"a5";
            when "00" & x"03c" => data <= x"b3";
            when "00" & x"03d" => data <= x"48";
            when "00" & x"03e" => data <= x"98";
            when "00" & x"03f" => data <= x"48";
            when "00" & x"040" => data <= x"a0";
            when "00" & x"041" => data <= x"00";
            when "00" & x"042" => data <= x"20";
            when "00" & x"043" => data <= x"da";
            when "00" & x"044" => data <= x"83";
            when "00" & x"045" => data <= x"b1";
            when "00" & x"046" => data <= x"ae";
            when "00" & x"047" => data <= x"8d";
            when "00" & x"048" => data <= x"01";
            when "00" & x"049" => data <= x"01";
            when "00" & x"04a" => data <= x"2c";
            when "00" & x"04b" => data <= x"de";
            when "00" & x"04c" => data <= x"10";
            when "00" & x"04d" => data <= x"10";
            when "00" & x"04e" => data <= x"25";
            when "00" & x"04f" => data <= x"a9";
            when "00" & x"050" => data <= x"02";
            when "00" & x"051" => data <= x"8d";
            when "00" & x"052" => data <= x"de";
            when "00" & x"053" => data <= x"10";
            when "00" & x"054" => data <= x"a9";
            when "00" & x"055" => data <= x"00";
            when "00" & x"056" => data <= x"8d";
            when "00" & x"057" => data <= x"00";
            when "00" & x"058" => data <= x"01";
            when "00" & x"059" => data <= x"f0";
            when "00" & x"05a" => data <= x"19";
            when "00" & x"05b" => data <= x"a9";
            when "00" & x"05c" => data <= x"02";
            when "00" & x"05d" => data <= x"8d";
            when "00" & x"05e" => data <= x"de";
            when "00" & x"05f" => data <= x"10";
            when "00" & x"060" => data <= x"a9";
            when "00" & x"061" => data <= x"00";
            when "00" & x"062" => data <= x"8d";
            when "00" & x"063" => data <= x"00";
            when "00" & x"064" => data <= x"01";
            when "00" & x"065" => data <= x"85";
            when "00" & x"066" => data <= x"b3";
            when "00" & x"067" => data <= x"68";
            when "00" & x"068" => data <= x"85";
            when "00" & x"069" => data <= x"ae";
            when "00" & x"06a" => data <= x"68";
            when "00" & x"06b" => data <= x"85";
            when "00" & x"06c" => data <= x"af";
            when "00" & x"06d" => data <= x"a5";
            when "00" & x"06e" => data <= x"b3";
            when "00" & x"06f" => data <= x"48";
            when "00" & x"070" => data <= x"98";
            when "00" & x"071" => data <= x"48";
            when "00" & x"072" => data <= x"a0";
            when "00" & x"073" => data <= x"00";
            when "00" & x"074" => data <= x"20";
            when "00" & x"075" => data <= x"da";
            when "00" & x"076" => data <= x"83";
            when "00" & x"077" => data <= x"b1";
            when "00" & x"078" => data <= x"ae";
            when "00" & x"079" => data <= x"30";
            when "00" & x"07a" => data <= x"08";
            when "00" & x"07b" => data <= x"f0";
            when "00" & x"07c" => data <= x"0d";
            when "00" & x"07d" => data <= x"20";
            when "00" & x"07e" => data <= x"9c";
            when "00" & x"07f" => data <= x"80";
            when "00" & x"080" => data <= x"4c";
            when "00" & x"081" => data <= x"74";
            when "00" & x"082" => data <= x"80";
            when "00" & x"083" => data <= x"68";
            when "00" & x"084" => data <= x"a8";
            when "00" & x"085" => data <= x"68";
            when "00" & x"086" => data <= x"18";
            when "00" & x"087" => data <= x"6c";
            when "00" & x"088" => data <= x"ae";
            when "00" & x"089" => data <= x"00";
            when "00" & x"08a" => data <= x"a9";
            when "00" & x"08b" => data <= x"00";
            when "00" & x"08c" => data <= x"ae";
            when "00" & x"08d" => data <= x"de";
            when "00" & x"08e" => data <= x"10";
            when "00" & x"08f" => data <= x"9d";
            when "00" & x"090" => data <= x"00";
            when "00" & x"091" => data <= x"01";
            when "00" & x"092" => data <= x"a9";
            when "00" & x"093" => data <= x"ff";
            when "00" & x"094" => data <= x"8d";
            when "00" & x"095" => data <= x"de";
            when "00" & x"096" => data <= x"10";
            when "00" & x"097" => data <= x"4c";
            when "00" & x"098" => data <= x"00";
            when "00" & x"099" => data <= x"01";
            when "00" & x"09a" => data <= x"a9";
            when "00" & x"09b" => data <= x"2e";
            when "00" & x"09c" => data <= x"20";
            when "00" & x"09d" => data <= x"e1";
            when "00" & x"09e" => data <= x"83";
            when "00" & x"09f" => data <= x"2c";
            when "00" & x"0a0" => data <= x"de";
            when "00" & x"0a1" => data <= x"10";
            when "00" & x"0a2" => data <= x"10";
            when "00" & x"0a3" => data <= x"14";
            when "00" & x"0a4" => data <= x"48";
            when "00" & x"0a5" => data <= x"20";
            when "00" & x"0a6" => data <= x"1c";
            when "00" & x"0a7" => data <= x"99";
            when "00" & x"0a8" => data <= x"8a";
            when "00" & x"0a9" => data <= x"48";
            when "00" & x"0aa" => data <= x"09";
            when "00" & x"0ab" => data <= x"10";
            when "00" & x"0ac" => data <= x"20";
            when "00" & x"0ad" => data <= x"17";
            when "00" & x"0ae" => data <= x"99";
            when "00" & x"0af" => data <= x"68";
            when "00" & x"0b0" => data <= x"aa";
            when "00" & x"0b1" => data <= x"68";
            when "00" & x"0b2" => data <= x"20";
            when "00" & x"0b3" => data <= x"e3";
            when "00" & x"0b4" => data <= x"ff";
            when "00" & x"0b5" => data <= x"4c";
            when "00" & x"0b6" => data <= x"18";
            when "00" & x"0b7" => data <= x"99";
            when "00" & x"0b8" => data <= x"ae";
            when "00" & x"0b9" => data <= x"de";
            when "00" & x"0ba" => data <= x"10";
            when "00" & x"0bb" => data <= x"9d";
            when "00" & x"0bc" => data <= x"00";
            when "00" & x"0bd" => data <= x"01";
            when "00" & x"0be" => data <= x"ee";
            when "00" & x"0bf" => data <= x"de";
            when "00" & x"0c0" => data <= x"10";
            when "00" & x"0c1" => data <= x"60";
            when "00" & x"0c2" => data <= x"48";
            when "00" & x"0c3" => data <= x"20";
            when "00" & x"0c4" => data <= x"05";
            when "00" & x"0c5" => data <= x"82";
            when "00" & x"0c6" => data <= x"20";
            when "00" & x"0c7" => data <= x"ca";
            when "00" & x"0c8" => data <= x"80";
            when "00" & x"0c9" => data <= x"68";
            when "00" & x"0ca" => data <= x"48";
            when "00" & x"0cb" => data <= x"29";
            when "00" & x"0cc" => data <= x"0f";
            when "00" & x"0cd" => data <= x"c9";
            when "00" & x"0ce" => data <= x"0a";
            when "00" & x"0cf" => data <= x"90";
            when "00" & x"0d0" => data <= x"02";
            when "00" & x"0d1" => data <= x"69";
            when "00" & x"0d2" => data <= x"06";
            when "00" & x"0d3" => data <= x"69";
            when "00" & x"0d4" => data <= x"30";
            when "00" & x"0d5" => data <= x"20";
            when "00" & x"0d6" => data <= x"9c";
            when "00" & x"0d7" => data <= x"80";
            when "00" & x"0d8" => data <= x"68";
            when "00" & x"0d9" => data <= x"60";
            when "00" & x"0da" => data <= x"20";
            when "00" & x"0db" => data <= x"ea";
            when "00" & x"0dc" => data <= x"80";
            when "00" & x"0dd" => data <= x"ca";
            when "00" & x"0de" => data <= x"ca";
            when "00" & x"0df" => data <= x"20";
            when "00" & x"0e0" => data <= x"e2";
            when "00" & x"0e1" => data <= x"80";
            when "00" & x"0e2" => data <= x"b1";
            when "00" & x"0e3" => data <= x"b0";
            when "00" & x"0e4" => data <= x"9d";
            when "00" & x"0e5" => data <= x"72";
            when "00" & x"0e6" => data <= x"10";
            when "00" & x"0e7" => data <= x"e8";
            when "00" & x"0e8" => data <= x"c8";
            when "00" & x"0e9" => data <= x"60";
            when "00" & x"0ea" => data <= x"20";
            when "00" & x"0eb" => data <= x"ed";
            when "00" & x"0ec" => data <= x"80";
            when "00" & x"0ed" => data <= x"b1";
            when "00" & x"0ee" => data <= x"b0";
            when "00" & x"0ef" => data <= x"95";
            when "00" & x"0f0" => data <= x"bc";
            when "00" & x"0f1" => data <= x"e8";
            when "00" & x"0f2" => data <= x"c8";
            when "00" & x"0f3" => data <= x"60";
            when "00" & x"0f4" => data <= x"a9";
            when "00" & x"0f5" => data <= x"20";
            when "00" & x"0f6" => data <= x"a2";
            when "00" & x"0f7" => data <= x"06";
            when "00" & x"0f8" => data <= x"95";
            when "00" & x"0f9" => data <= x"c7";
            when "00" & x"0fa" => data <= x"ca";
            when "00" & x"0fb" => data <= x"10";
            when "00" & x"0fc" => data <= x"fb";
            when "00" & x"0fd" => data <= x"60";
            when "00" & x"0fe" => data <= x"20";
            when "00" & x"0ff" => data <= x"4d";
            when "00" & x"100" => data <= x"83";
            when "00" & x"101" => data <= x"20";
            when "00" & x"102" => data <= x"f4";
            when "00" & x"103" => data <= x"80";
            when "00" & x"104" => data <= x"30";
            when "00" & x"105" => data <= x"13";
            when "00" & x"106" => data <= x"20";
            when "00" & x"107" => data <= x"4d";
            when "00" & x"108" => data <= x"83";
            when "00" & x"109" => data <= x"20";
            when "00" & x"10a" => data <= x"f4";
            when "00" & x"10b" => data <= x"80";
            when "00" & x"10c" => data <= x"a5";
            when "00" & x"10d" => data <= x"bc";
            when "00" & x"10e" => data <= x"85";
            when "00" & x"10f" => data <= x"f2";
            when "00" & x"110" => data <= x"a5";
            when "00" & x"111" => data <= x"bd";
            when "00" & x"112" => data <= x"85";
            when "00" & x"113" => data <= x"f3";
            when "00" & x"114" => data <= x"a0";
            when "00" & x"115" => data <= x"00";
            when "00" & x"116" => data <= x"20";
            when "00" & x"117" => data <= x"bf";
            when "00" & x"118" => data <= x"86";
            when "00" & x"119" => data <= x"a2";
            when "00" & x"11a" => data <= x"01";
            when "00" & x"11b" => data <= x"20";
            when "00" & x"11c" => data <= x"c5";
            when "00" & x"11d" => data <= x"ff";
            when "00" & x"11e" => data <= x"b0";
            when "00" & x"11f" => data <= x"dd";
            when "00" & x"120" => data <= x"85";
            when "00" & x"121" => data <= x"c7";
            when "00" & x"122" => data <= x"c9";
            when "00" & x"123" => data <= x"2e";
            when "00" & x"124" => data <= x"d0";
            when "00" & x"125" => data <= x"04";
            when "00" & x"126" => data <= x"a9";
            when "00" & x"127" => data <= x"20";
            when "00" & x"128" => data <= x"d0";
            when "00" & x"129" => data <= x"4d";
            when "00" & x"12a" => data <= x"c9";
            when "00" & x"12b" => data <= x"3a";
            when "00" & x"12c" => data <= x"d0";
            when "00" & x"12d" => data <= x"21";
            when "00" & x"12e" => data <= x"20";
            when "00" & x"12f" => data <= x"c5";
            when "00" & x"130" => data <= x"ff";
            when "00" & x"131" => data <= x"b0";
            when "00" & x"132" => data <= x"15";
            when "00" & x"133" => data <= x"38";
            when "00" & x"134" => data <= x"e9";
            when "00" & x"135" => data <= x"30";
            when "00" & x"136" => data <= x"90";
            when "00" & x"137" => data <= x"10";
            when "00" & x"138" => data <= x"c9";
            when "00" & x"139" => data <= x"04";
            when "00" & x"13a" => data <= x"b0";
            when "00" & x"13b" => data <= x"0c";
            when "00" & x"13c" => data <= x"20";
            when "00" & x"13d" => data <= x"7e";
            when "00" & x"13e" => data <= x"87";
            when "00" & x"13f" => data <= x"20";
            when "00" & x"140" => data <= x"c5";
            when "00" & x"141" => data <= x"ff";
            when "00" & x"142" => data <= x"b0";
            when "00" & x"143" => data <= x"5c";
            when "00" & x"144" => data <= x"c9";
            when "00" & x"145" => data <= x"2e";
            when "00" & x"146" => data <= x"f0";
            when "00" & x"147" => data <= x"03";
            when "00" & x"148" => data <= x"4c";
            when "00" & x"149" => data <= x"74";
            when "00" & x"14a" => data <= x"83";
            when "00" & x"14b" => data <= x"a9";
            when "00" & x"14c" => data <= x"24";
            when "00" & x"14d" => data <= x"d0";
            when "00" & x"14e" => data <= x"28";
            when "00" & x"14f" => data <= x"c9";
            when "00" & x"150" => data <= x"2a";
            when "00" & x"151" => data <= x"d0";
            when "00" & x"152" => data <= x"19";
            when "00" & x"153" => data <= x"20";
            when "00" & x"154" => data <= x"c5";
            when "00" & x"155" => data <= x"ff";
            when "00" & x"156" => data <= x"b0";
            when "00" & x"157" => data <= x"08";
            when "00" & x"158" => data <= x"c9";
            when "00" & x"159" => data <= x"2e";
            when "00" & x"15a" => data <= x"d0";
            when "00" & x"15b" => data <= x"32";
            when "00" & x"15c" => data <= x"a9";
            when "00" & x"15d" => data <= x"23";
            when "00" & x"15e" => data <= x"d0";
            when "00" & x"15f" => data <= x"17";
            when "00" & x"160" => data <= x"a2";
            when "00" & x"161" => data <= x"00";
            when "00" & x"162" => data <= x"a9";
            when "00" & x"163" => data <= x"23";
            when "00" & x"164" => data <= x"95";
            when "00" & x"165" => data <= x"c7";
            when "00" & x"166" => data <= x"e8";
            when "00" & x"167" => data <= x"e0";
            when "00" & x"168" => data <= x"07";
            when "00" & x"169" => data <= x"d0";
            when "00" & x"16a" => data <= x"f9";
            when "00" & x"16b" => data <= x"60";
            when "00" & x"16c" => data <= x"20";
            when "00" & x"16d" => data <= x"c5";
            when "00" & x"16e" => data <= x"ff";
            when "00" & x"16f" => data <= x"b0";
            when "00" & x"170" => data <= x"2f";
            when "00" & x"171" => data <= x"c9";
            when "00" & x"172" => data <= x"2e";
            when "00" & x"173" => data <= x"d0";
            when "00" & x"174" => data <= x"10";
            when "00" & x"175" => data <= x"a5";
            when "00" & x"176" => data <= x"c7";
            when "00" & x"177" => data <= x"85";
            when "00" & x"178" => data <= x"ce";
            when "00" & x"179" => data <= x"4c";
            when "00" & x"17a" => data <= x"1b";
            when "00" & x"17b" => data <= x"81";
            when "00" & x"17c" => data <= x"20";
            when "00" & x"17d" => data <= x"c5";
            when "00" & x"17e" => data <= x"ff";
            when "00" & x"17f" => data <= x"b0";
            when "00" & x"180" => data <= x"1f";
            when "00" & x"181" => data <= x"e0";
            when "00" & x"182" => data <= x"07";
            when "00" & x"183" => data <= x"f0";
            when "00" & x"184" => data <= x"09";
            when "00" & x"185" => data <= x"c9";
            when "00" & x"186" => data <= x"2a";
            when "00" & x"187" => data <= x"d0";
            when "00" & x"188" => data <= x"12";
            when "00" & x"189" => data <= x"20";
            when "00" & x"18a" => data <= x"c5";
            when "00" & x"18b" => data <= x"ff";
            when "00" & x"18c" => data <= x"b0";
            when "00" & x"18d" => data <= x"d4";
            when "00" & x"18e" => data <= x"20";
            when "00" & x"18f" => data <= x"22";
            when "00" & x"190" => data <= x"80";
            when "00" & x"191" => data <= x"cc";
            when "00" & x"192" => data <= x"66";
            when "00" & x"193" => data <= x"69";
            when "00" & x"194" => data <= x"6c";
            when "00" & x"195" => data <= x"65";
            when "00" & x"196" => data <= x"6e";
            when "00" & x"197" => data <= x"61";
            when "00" & x"198" => data <= x"6d";
            when "00" & x"199" => data <= x"65";
            when "00" & x"19a" => data <= x"00";
            when "00" & x"19b" => data <= x"95";
            when "00" & x"19c" => data <= x"c7";
            when "00" & x"19d" => data <= x"e8";
            when "00" & x"19e" => data <= x"d0";
            when "00" & x"19f" => data <= x"dc";
            when "00" & x"1a0" => data <= x"60";
            when "00" & x"1a1" => data <= x"20";
            when "00" & x"1a2" => data <= x"e1";
            when "00" & x"1a3" => data <= x"83";
            when "00" & x"1a4" => data <= x"ad";
            when "00" & x"1a5" => data <= x"04";
            when "00" & x"1a6" => data <= x"0f";
            when "00" & x"1a7" => data <= x"20";
            when "00" & x"1a8" => data <= x"47";
            when "00" & x"1a9" => data <= x"83";
            when "00" & x"1aa" => data <= x"cd";
            when "00" & x"1ab" => data <= x"04";
            when "00" & x"1ac" => data <= x"0f";
            when "00" & x"1ad" => data <= x"f0";
            when "00" & x"1ae" => data <= x"f1";
            when "00" & x"1af" => data <= x"20";
            when "00" & x"1b0" => data <= x"33";
            when "00" & x"1b1" => data <= x"80";
            when "00" & x"1b2" => data <= x"c8";
            when "00" & x"1b3" => data <= x"44";
            when "00" & x"1b4" => data <= x"69";
            when "00" & x"1b5" => data <= x"73";
            when "00" & x"1b6" => data <= x"6b";
            when "00" & x"1b7" => data <= x"20";
            when "00" & x"1b8" => data <= x"63";
            when "00" & x"1b9" => data <= x"68";
            when "00" & x"1ba" => data <= x"61";
            when "00" & x"1bb" => data <= x"6e";
            when "00" & x"1bc" => data <= x"67";
            when "00" & x"1bd" => data <= x"65";
            when "00" & x"1be" => data <= x"64";
            when "00" & x"1bf" => data <= x"00";
            when "00" & x"1c0" => data <= x"20";
            when "00" & x"1c1" => data <= x"e1";
            when "00" & x"1c2" => data <= x"83";
            when "00" & x"1c3" => data <= x"b9";
            when "00" & x"1c4" => data <= x"0f";
            when "00" & x"1c5" => data <= x"0e";
            when "00" & x"1c6" => data <= x"08";
            when "00" & x"1c7" => data <= x"29";
            when "00" & x"1c8" => data <= x"7f";
            when "00" & x"1c9" => data <= x"d0";
            when "00" & x"1ca" => data <= x"05";
            when "00" & x"1cb" => data <= x"20";
            when "00" & x"1cc" => data <= x"cb";
            when "00" & x"1cd" => data <= x"9f";
            when "00" & x"1ce" => data <= x"f0";
            when "00" & x"1cf" => data <= x"06";
            when "00" & x"1d0" => data <= x"20";
            when "00" & x"1d1" => data <= x"9c";
            when "00" & x"1d2" => data <= x"80";
            when "00" & x"1d3" => data <= x"20";
            when "00" & x"1d4" => data <= x"9a";
            when "00" & x"1d5" => data <= x"80";
            when "00" & x"1d6" => data <= x"a2";
            when "00" & x"1d7" => data <= x"06";
            when "00" & x"1d8" => data <= x"b9";
            when "00" & x"1d9" => data <= x"08";
            when "00" & x"1da" => data <= x"0e";
            when "00" & x"1db" => data <= x"29";
            when "00" & x"1dc" => data <= x"7f";
            when "00" & x"1dd" => data <= x"20";
            when "00" & x"1de" => data <= x"9c";
            when "00" & x"1df" => data <= x"80";
            when "00" & x"1e0" => data <= x"c8";
            when "00" & x"1e1" => data <= x"ca";
            when "00" & x"1e2" => data <= x"10";
            when "00" & x"1e3" => data <= x"f4";
            when "00" & x"1e4" => data <= x"20";
            when "00" & x"1e5" => data <= x"cb";
            when "00" & x"1e6" => data <= x"9f";
            when "00" & x"1e7" => data <= x"a9";
            when "00" & x"1e8" => data <= x"20";
            when "00" & x"1e9" => data <= x"28";
            when "00" & x"1ea" => data <= x"10";
            when "00" & x"1eb" => data <= x"02";
            when "00" & x"1ec" => data <= x"a9";
            when "00" & x"1ed" => data <= x"4c";
            when "00" & x"1ee" => data <= x"20";
            when "00" & x"1ef" => data <= x"9c";
            when "00" & x"1f0" => data <= x"80";
            when "00" & x"1f1" => data <= x"4c";
            when "00" & x"1f2" => data <= x"ce";
            when "00" & x"1f3" => data <= x"9f";
            when "00" & x"1f4" => data <= x"20";
            when "00" & x"1f5" => data <= x"ce";
            when "00" & x"1f6" => data <= x"9f";
            when "00" & x"1f7" => data <= x"88";
            when "00" & x"1f8" => data <= x"d0";
            when "00" & x"1f9" => data <= x"fa";
            when "00" & x"1fa" => data <= x"60";
            when "00" & x"1fb" => data <= x"4a";
            when "00" & x"1fc" => data <= x"4a";
            when "00" & x"1fd" => data <= x"4a";
            when "00" & x"1fe" => data <= x"4a";
            when "00" & x"1ff" => data <= x"4a";
            when "00" & x"200" => data <= x"4a";
            when "00" & x"201" => data <= x"29";
            when "00" & x"202" => data <= x"03";
            when "00" & x"203" => data <= x"60";
            when "00" & x"204" => data <= x"4a";
            when "00" & x"205" => data <= x"4a";
            when "00" & x"206" => data <= x"4a";
            when "00" & x"207" => data <= x"4a";
            when "00" & x"208" => data <= x"4a";
            when "00" & x"209" => data <= x"60";
            when "00" & x"20a" => data <= x"0a";
            when "00" & x"20b" => data <= x"0a";
            when "00" & x"20c" => data <= x"0a";
            when "00" & x"20d" => data <= x"0a";
            when "00" & x"20e" => data <= x"0a";
            when "00" & x"20f" => data <= x"60";
            when "00" & x"210" => data <= x"c8";
            when "00" & x"211" => data <= x"c8";
            when "00" & x"212" => data <= x"c8";
            when "00" & x"213" => data <= x"c8";
            when "00" & x"214" => data <= x"c8";
            when "00" & x"215" => data <= x"c8";
            when "00" & x"216" => data <= x"c8";
            when "00" & x"217" => data <= x"c8";
            when "00" & x"218" => data <= x"60";
            when "00" & x"219" => data <= x"88";
            when "00" & x"21a" => data <= x"88";
            when "00" & x"21b" => data <= x"88";
            when "00" & x"21c" => data <= x"88";
            when "00" & x"21d" => data <= x"88";
            when "00" & x"21e" => data <= x"88";
            when "00" & x"21f" => data <= x"88";
            when "00" & x"220" => data <= x"88";
            when "00" & x"221" => data <= x"60";
            when "00" & x"222" => data <= x"00";
            when "00" & x"223" => data <= x"00";
            when "00" & x"224" => data <= x"00";
            when "00" & x"225" => data <= x"00";
            when "00" & x"226" => data <= x"00";
            when "00" & x"227" => data <= x"00";
            when "00" & x"228" => data <= x"00";
            when "00" & x"229" => data <= x"00";
            when "00" & x"22a" => data <= x"00";
            when "00" & x"22b" => data <= x"00";
            when "00" & x"22c" => data <= x"00";
            when "00" & x"22d" => data <= x"00";
            when "00" & x"22e" => data <= x"00";
            when "00" & x"22f" => data <= x"00";
            when "00" & x"230" => data <= x"00";
            when "00" & x"231" => data <= x"00";
            when "00" & x"232" => data <= x"00";
            when "00" & x"233" => data <= x"00";
            when "00" & x"234" => data <= x"00";
            when "00" & x"235" => data <= x"00";
            when "00" & x"236" => data <= x"00";
            when "00" & x"237" => data <= x"00";
            when "00" & x"238" => data <= x"00";
            when "00" & x"239" => data <= x"00";
            when "00" & x"23a" => data <= x"00";
            when "00" & x"23b" => data <= x"00";
            when "00" & x"23c" => data <= x"00";
            when "00" & x"23d" => data <= x"00";
            when "00" & x"23e" => data <= x"00";
            when "00" & x"23f" => data <= x"00";
            when "00" & x"240" => data <= x"00";
            when "00" & x"241" => data <= x"00";
            when "00" & x"242" => data <= x"00";
            when "00" & x"243" => data <= x"00";
            when "00" & x"244" => data <= x"00";
            when "00" & x"245" => data <= x"00";
            when "00" & x"246" => data <= x"00";
            when "00" & x"247" => data <= x"00";
            when "00" & x"248" => data <= x"00";
            when "00" & x"249" => data <= x"00";
            when "00" & x"24a" => data <= x"00";
            when "00" & x"24b" => data <= x"00";
            when "00" & x"24c" => data <= x"00";
            when "00" & x"24d" => data <= x"00";
            when "00" & x"24e" => data <= x"00";
            when "00" & x"24f" => data <= x"00";
            when "00" & x"250" => data <= x"00";
            when "00" & x"251" => data <= x"00";
            when "00" & x"252" => data <= x"00";
            when "00" & x"253" => data <= x"00";
            when "00" & x"254" => data <= x"00";
            when "00" & x"255" => data <= x"00";
            when "00" & x"256" => data <= x"00";
            when "00" & x"257" => data <= x"00";
            when "00" & x"258" => data <= x"00";
            when "00" & x"259" => data <= x"00";
            when "00" & x"25a" => data <= x"00";
            when "00" & x"25b" => data <= x"00";
            when "00" & x"25c" => data <= x"00";
            when "00" & x"25d" => data <= x"60";
            when "00" & x"25e" => data <= x"a9";
            when "00" & x"25f" => data <= x"23";
            when "00" & x"260" => data <= x"d0";
            when "00" & x"261" => data <= x"02";
            when "00" & x"262" => data <= x"a9";
            when "00" & x"263" => data <= x"ff";
            when "00" & x"264" => data <= x"8d";
            when "00" & x"265" => data <= x"cf";
            when "00" & x"266" => data <= x"10";
            when "00" & x"267" => data <= x"60";
            when "00" & x"268" => data <= x"20";
            when "00" & x"269" => data <= x"fe";
            when "00" & x"26a" => data <= x"80";
            when "00" & x"26b" => data <= x"4c";
            when "00" & x"26c" => data <= x"71";
            when "00" & x"26d" => data <= x"82";
            when "00" & x"26e" => data <= x"20";
            when "00" & x"26f" => data <= x"06";
            when "00" & x"270" => data <= x"81";
            when "00" & x"271" => data <= x"20";
            when "00" & x"272" => data <= x"96";
            when "00" & x"273" => data <= x"82";
            when "00" & x"274" => data <= x"b0";
            when "00" & x"275" => data <= x"e7";
            when "00" & x"276" => data <= x"20";
            when "00" & x"277" => data <= x"2b";
            when "00" & x"278" => data <= x"80";
            when "00" & x"279" => data <= x"d6";
            when "00" & x"27a" => data <= x"6e";
            when "00" & x"27b" => data <= x"6f";
            when "00" & x"27c" => data <= x"74";
            when "00" & x"27d" => data <= x"20";
            when "00" & x"27e" => data <= x"66";
            when "00" & x"27f" => data <= x"6f";
            when "00" & x"280" => data <= x"75";
            when "00" & x"281" => data <= x"6e";
            when "00" & x"282" => data <= x"64";
            when "00" & x"283" => data <= x"00";
            when "00" & x"284" => data <= x"20";
            when "00" & x"285" => data <= x"5e";
            when "00" & x"286" => data <= x"82";
            when "00" & x"287" => data <= x"20";
            when "00" & x"288" => data <= x"01";
            when "00" & x"289" => data <= x"9a";
            when "00" & x"28a" => data <= x"20";
            when "00" & x"28b" => data <= x"68";
            when "00" & x"28c" => data <= x"82";
            when "00" & x"28d" => data <= x"20";
            when "00" & x"28e" => data <= x"01";
            when "00" & x"28f" => data <= x"83";
            when "00" & x"290" => data <= x"20";
            when "00" & x"291" => data <= x"9d";
            when "00" & x"292" => data <= x"82";
            when "00" & x"293" => data <= x"b0";
            when "00" & x"294" => data <= x"f8";
            when "00" & x"295" => data <= x"60";
            when "00" & x"296" => data <= x"20";
            when "00" & x"297" => data <= x"41";
            when "00" & x"298" => data <= x"af";
            when "00" & x"299" => data <= x"a0";
            when "00" & x"29a" => data <= x"f8";
            when "00" & x"29b" => data <= x"d0";
            when "00" & x"29c" => data <= x"03";
            when "00" & x"29d" => data <= x"ac";
            when "00" & x"29e" => data <= x"ce";
            when "00" & x"29f" => data <= x"10";
            when "00" & x"2a0" => data <= x"20";
            when "00" & x"2a1" => data <= x"10";
            when "00" & x"2a2" => data <= x"82";
            when "00" & x"2a3" => data <= x"cc";
            when "00" & x"2a4" => data <= x"05";
            when "00" & x"2a5" => data <= x"0f";
            when "00" & x"2a6" => data <= x"b0";
            when "00" & x"2a7" => data <= x"44";
            when "00" & x"2a8" => data <= x"20";
            when "00" & x"2a9" => data <= x"10";
            when "00" & x"2aa" => data <= x"82";
            when "00" & x"2ab" => data <= x"a2";
            when "00" & x"2ac" => data <= x"07";
            when "00" & x"2ad" => data <= x"b5";
            when "00" & x"2ae" => data <= x"c7";
            when "00" & x"2af" => data <= x"cd";
            when "00" & x"2b0" => data <= x"cf";
            when "00" & x"2b1" => data <= x"10";
            when "00" & x"2b2" => data <= x"f0";
            when "00" & x"2b3" => data <= x"0e";
            when "00" & x"2b4" => data <= x"20";
            when "00" & x"2b5" => data <= x"ee";
            when "00" & x"2b6" => data <= x"82";
            when "00" & x"2b7" => data <= x"59";
            when "00" & x"2b8" => data <= x"07";
            when "00" & x"2b9" => data <= x"0e";
            when "00" & x"2ba" => data <= x"b0";
            when "00" & x"2bb" => data <= x"02";
            when "00" & x"2bc" => data <= x"29";
            when "00" & x"2bd" => data <= x"df";
            when "00" & x"2be" => data <= x"29";
            when "00" & x"2bf" => data <= x"7f";
            when "00" & x"2c0" => data <= x"d0";
            when "00" & x"2c1" => data <= x"09";
            when "00" & x"2c2" => data <= x"88";
            when "00" & x"2c3" => data <= x"ca";
            when "00" & x"2c4" => data <= x"10";
            when "00" & x"2c5" => data <= x"e7";
            when "00" & x"2c6" => data <= x"8c";
            when "00" & x"2c7" => data <= x"ce";
            when "00" & x"2c8" => data <= x"10";
            when "00" & x"2c9" => data <= x"38";
            when "00" & x"2ca" => data <= x"60";
            when "00" & x"2cb" => data <= x"88";
            when "00" & x"2cc" => data <= x"ca";
            when "00" & x"2cd" => data <= x"10";
            when "00" & x"2ce" => data <= x"fc";
            when "00" & x"2cf" => data <= x"30";
            when "00" & x"2d0" => data <= x"cf";
            when "00" & x"2d1" => data <= x"20";
            when "00" & x"2d2" => data <= x"4c";
            when "00" & x"2d3" => data <= x"98";
            when "00" & x"2d4" => data <= x"b9";
            when "00" & x"2d5" => data <= x"10";
            when "00" & x"2d6" => data <= x"0e";
            when "00" & x"2d7" => data <= x"99";
            when "00" & x"2d8" => data <= x"08";
            when "00" & x"2d9" => data <= x"0e";
            when "00" & x"2da" => data <= x"b9";
            when "00" & x"2db" => data <= x"10";
            when "00" & x"2dc" => data <= x"0f";
            when "00" & x"2dd" => data <= x"99";
            when "00" & x"2de" => data <= x"08";
            when "00" & x"2df" => data <= x"0f";
            when "00" & x"2e0" => data <= x"c8";
            when "00" & x"2e1" => data <= x"cc";
            when "00" & x"2e2" => data <= x"05";
            when "00" & x"2e3" => data <= x"0f";
            when "00" & x"2e4" => data <= x"90";
            when "00" & x"2e5" => data <= x"ee";
            when "00" & x"2e6" => data <= x"98";
            when "00" & x"2e7" => data <= x"e9";
            when "00" & x"2e8" => data <= x"08";
            when "00" & x"2e9" => data <= x"8d";
            when "00" & x"2ea" => data <= x"05";
            when "00" & x"2eb" => data <= x"0f";
            when "00" & x"2ec" => data <= x"18";
            when "00" & x"2ed" => data <= x"60";
            when "00" & x"2ee" => data <= x"48";
            when "00" & x"2ef" => data <= x"29";
            when "00" & x"2f0" => data <= x"df";
            when "00" & x"2f1" => data <= x"c9";
            when "00" & x"2f2" => data <= x"41";
            when "00" & x"2f3" => data <= x"90";
            when "00" & x"2f4" => data <= x"04";
            when "00" & x"2f5" => data <= x"c9";
            when "00" & x"2f6" => data <= x"5b";
            when "00" & x"2f7" => data <= x"90";
            when "00" & x"2f8" => data <= x"01";
            when "00" & x"2f9" => data <= x"38";
            when "00" & x"2fa" => data <= x"68";
            when "00" & x"2fb" => data <= x"60";
            when "00" & x"2fc" => data <= x"2c";
            when "00" & x"2fd" => data <= x"c7";
            when "00" & x"2fe" => data <= x"10";
            when "00" & x"2ff" => data <= x"30";
            when "00" & x"300" => data <= x"ec";
            when "00" & x"301" => data <= x"20";
            when "00" & x"302" => data <= x"e1";
            when "00" & x"303" => data <= x"83";
            when "00" & x"304" => data <= x"20";
            when "00" & x"305" => data <= x"c0";
            when "00" & x"306" => data <= x"81";
            when "00" & x"307" => data <= x"98";
            when "00" & x"308" => data <= x"48";
            when "00" & x"309" => data <= x"a9";
            when "00" & x"30a" => data <= x"60";
            when "00" & x"30b" => data <= x"85";
            when "00" & x"30c" => data <= x"b0";
            when "00" & x"30d" => data <= x"a9";
            when "00" & x"30e" => data <= x"10";
            when "00" & x"30f" => data <= x"85";
            when "00" & x"310" => data <= x"b1";
            when "00" & x"311" => data <= x"20";
            when "00" & x"312" => data <= x"7e";
            when "00" & x"313" => data <= x"83";
            when "00" & x"314" => data <= x"a0";
            when "00" & x"315" => data <= x"02";
            when "00" & x"316" => data <= x"20";
            when "00" & x"317" => data <= x"ce";
            when "00" & x"318" => data <= x"9f";
            when "00" & x"319" => data <= x"20";
            when "00" & x"31a" => data <= x"35";
            when "00" & x"31b" => data <= x"83";
            when "00" & x"31c" => data <= x"20";
            when "00" & x"31d" => data <= x"35";
            when "00" & x"31e" => data <= x"83";
            when "00" & x"31f" => data <= x"20";
            when "00" & x"320" => data <= x"35";
            when "00" & x"321" => data <= x"83";
            when "00" & x"322" => data <= x"68";
            when "00" & x"323" => data <= x"a8";
            when "00" & x"324" => data <= x"b9";
            when "00" & x"325" => data <= x"0e";
            when "00" & x"326" => data <= x"0f";
            when "00" & x"327" => data <= x"29";
            when "00" & x"328" => data <= x"03";
            when "00" & x"329" => data <= x"20";
            when "00" & x"32a" => data <= x"ca";
            when "00" & x"32b" => data <= x"80";
            when "00" & x"32c" => data <= x"b9";
            when "00" & x"32d" => data <= x"0f";
            when "00" & x"32e" => data <= x"0f";
            when "00" & x"32f" => data <= x"20";
            when "00" & x"330" => data <= x"c2";
            when "00" & x"331" => data <= x"80";
            when "00" & x"332" => data <= x"4c";
            when "00" & x"333" => data <= x"9a";
            when "00" & x"334" => data <= x"9f";
            when "00" & x"335" => data <= x"a2";
            when "00" & x"336" => data <= x"03";
            when "00" & x"337" => data <= x"b9";
            when "00" & x"338" => data <= x"62";
            when "00" & x"339" => data <= x"10";
            when "00" & x"33a" => data <= x"20";
            when "00" & x"33b" => data <= x"c2";
            when "00" & x"33c" => data <= x"80";
            when "00" & x"33d" => data <= x"88";
            when "00" & x"33e" => data <= x"ca";
            when "00" & x"33f" => data <= x"d0";
            when "00" & x"340" => data <= x"f6";
            when "00" & x"341" => data <= x"20";
            when "00" & x"342" => data <= x"11";
            when "00" & x"343" => data <= x"82";
            when "00" & x"344" => data <= x"4c";
            when "00" & x"345" => data <= x"ce";
            when "00" & x"346" => data <= x"9f";
            when "00" & x"347" => data <= x"20";
            when "00" & x"348" => data <= x"e1";
            when "00" & x"349" => data <= x"83";
            when "00" & x"34a" => data <= x"4c";
            when "00" & x"34b" => data <= x"41";
            when "00" & x"34c" => data <= x"af";
            when "00" & x"34d" => data <= x"ad";
            when "00" & x"34e" => data <= x"ca";
            when "00" & x"34f" => data <= x"10";
            when "00" & x"350" => data <= x"85";
            when "00" & x"351" => data <= x"ce";
            when "00" & x"352" => data <= x"ad";
            when "00" & x"353" => data <= x"cb";
            when "00" & x"354" => data <= x"10";
            when "00" & x"355" => data <= x"4c";
            when "00" & x"356" => data <= x"7e";
            when "00" & x"357" => data <= x"87";
            when "00" & x"358" => data <= x"20";
            when "00" & x"359" => data <= x"bf";
            when "00" & x"35a" => data <= x"86";
            when "00" & x"35b" => data <= x"f0";
            when "00" & x"35c" => data <= x"f5";
            when "00" & x"35d" => data <= x"20";
            when "00" & x"35e" => data <= x"c5";
            when "00" & x"35f" => data <= x"ff";
            when "00" & x"360" => data <= x"b0";
            when "00" & x"361" => data <= x"12";
            when "00" & x"362" => data <= x"c9";
            when "00" & x"363" => data <= x"3a";
            when "00" & x"364" => data <= x"f0";
            when "00" & x"365" => data <= x"f7";
            when "00" & x"366" => data <= x"38";
            when "00" & x"367" => data <= x"e9";
            when "00" & x"368" => data <= x"30";
            when "00" & x"369" => data <= x"90";
            when "00" & x"36a" => data <= x"09";
            when "00" & x"36b" => data <= x"c9";
            when "00" & x"36c" => data <= x"04";
            when "00" & x"36d" => data <= x"b0";
            when "00" & x"36e" => data <= x"05";
            when "00" & x"36f" => data <= x"20";
            when "00" & x"370" => data <= x"7e";
            when "00" & x"371" => data <= x"87";
            when "00" & x"372" => data <= x"18";
            when "00" & x"373" => data <= x"60";
            when "00" & x"374" => data <= x"20";
            when "00" & x"375" => data <= x"22";
            when "00" & x"376" => data <= x"80";
            when "00" & x"377" => data <= x"cd";
            when "00" & x"378" => data <= x"64";
            when "00" & x"379" => data <= x"72";
            when "00" & x"37a" => data <= x"69";
            when "00" & x"37b" => data <= x"76";
            when "00" & x"37c" => data <= x"65";
            when "00" & x"37d" => data <= x"00";
            when "00" & x"37e" => data <= x"20";
            when "00" & x"37f" => data <= x"e1";
            when "00" & x"380" => data <= x"83";
            when "00" & x"381" => data <= x"98";
            when "00" & x"382" => data <= x"48";
            when "00" & x"383" => data <= x"aa";
            when "00" & x"384" => data <= x"a0";
            when "00" & x"385" => data <= x"02";
            when "00" & x"386" => data <= x"a9";
            when "00" & x"387" => data <= x"00";
            when "00" & x"388" => data <= x"91";
            when "00" & x"389" => data <= x"b0";
            when "00" & x"38a" => data <= x"c8";
            when "00" & x"38b" => data <= x"c0";
            when "00" & x"38c" => data <= x"12";
            when "00" & x"38d" => data <= x"d0";
            when "00" & x"38e" => data <= x"f9";
            when "00" & x"38f" => data <= x"a0";
            when "00" & x"390" => data <= x"02";
            when "00" & x"391" => data <= x"20";
            when "00" & x"392" => data <= x"cf";
            when "00" & x"393" => data <= x"83";
            when "00" & x"394" => data <= x"c8";
            when "00" & x"395" => data <= x"c8";
            when "00" & x"396" => data <= x"c0";
            when "00" & x"397" => data <= x"0e";
            when "00" & x"398" => data <= x"d0";
            when "00" & x"399" => data <= x"f7";
            when "00" & x"39a" => data <= x"68";
            when "00" & x"39b" => data <= x"aa";
            when "00" & x"39c" => data <= x"bd";
            when "00" & x"39d" => data <= x"0f";
            when "00" & x"39e" => data <= x"0e";
            when "00" & x"39f" => data <= x"10";
            when "00" & x"3a0" => data <= x"06";
            when "00" & x"3a1" => data <= x"a9";
            when "00" & x"3a2" => data <= x"0a";
            when "00" & x"3a3" => data <= x"a0";
            when "00" & x"3a4" => data <= x"0e";
            when "00" & x"3a5" => data <= x"91";
            when "00" & x"3a6" => data <= x"b0";
            when "00" & x"3a7" => data <= x"bd";
            when "00" & x"3a8" => data <= x"0e";
            when "00" & x"3a9" => data <= x"0f";
            when "00" & x"3aa" => data <= x"a0";
            when "00" & x"3ab" => data <= x"04";
            when "00" & x"3ac" => data <= x"20";
            when "00" & x"3ad" => data <= x"bb";
            when "00" & x"3ae" => data <= x"83";
            when "00" & x"3af" => data <= x"a0";
            when "00" & x"3b0" => data <= x"0c";
            when "00" & x"3b1" => data <= x"4a";
            when "00" & x"3b2" => data <= x"4a";
            when "00" & x"3b3" => data <= x"48";
            when "00" & x"3b4" => data <= x"29";
            when "00" & x"3b5" => data <= x"03";
            when "00" & x"3b6" => data <= x"91";
            when "00" & x"3b7" => data <= x"b0";
            when "00" & x"3b8" => data <= x"68";
            when "00" & x"3b9" => data <= x"a0";
            when "00" & x"3ba" => data <= x"08";
            when "00" & x"3bb" => data <= x"4a";
            when "00" & x"3bc" => data <= x"4a";
            when "00" & x"3bd" => data <= x"48";
            when "00" & x"3be" => data <= x"29";
            when "00" & x"3bf" => data <= x"03";
            when "00" & x"3c0" => data <= x"91";
            when "00" & x"3c1" => data <= x"b0";
            when "00" & x"3c2" => data <= x"c9";
            when "00" & x"3c3" => data <= x"03";
            when "00" & x"3c4" => data <= x"d0";
            when "00" & x"3c5" => data <= x"07";
            when "00" & x"3c6" => data <= x"a9";
            when "00" & x"3c7" => data <= x"ff";
            when "00" & x"3c8" => data <= x"91";
            when "00" & x"3c9" => data <= x"b0";
            when "00" & x"3ca" => data <= x"c8";
            when "00" & x"3cb" => data <= x"91";
            when "00" & x"3cc" => data <= x"b0";
            when "00" & x"3cd" => data <= x"68";
            when "00" & x"3ce" => data <= x"60";
            when "00" & x"3cf" => data <= x"20";
            when "00" & x"3d0" => data <= x"d2";
            when "00" & x"3d1" => data <= x"83";
            when "00" & x"3d2" => data <= x"bd";
            when "00" & x"3d3" => data <= x"08";
            when "00" & x"3d4" => data <= x"0f";
            when "00" & x"3d5" => data <= x"91";
            when "00" & x"3d6" => data <= x"b0";
            when "00" & x"3d7" => data <= x"e8";
            when "00" & x"3d8" => data <= x"c8";
            when "00" & x"3d9" => data <= x"60";
            when "00" & x"3da" => data <= x"e6";
            when "00" & x"3db" => data <= x"ae";
            when "00" & x"3dc" => data <= x"d0";
            when "00" & x"3dd" => data <= x"02";
            when "00" & x"3de" => data <= x"e6";
            when "00" & x"3df" => data <= x"af";
            when "00" & x"3e0" => data <= x"60";
            when "00" & x"3e1" => data <= x"48";
            when "00" & x"3e2" => data <= x"8a";
            when "00" & x"3e3" => data <= x"48";
            when "00" & x"3e4" => data <= x"98";
            when "00" & x"3e5" => data <= x"48";
            when "00" & x"3e6" => data <= x"a9";
            when "00" & x"3e7" => data <= x"84";
            when "00" & x"3e8" => data <= x"48";
            when "00" & x"3e9" => data <= x"a9";
            when "00" & x"3ea" => data <= x"03";
            when "00" & x"3eb" => data <= x"48";
            when "00" & x"3ec" => data <= x"a0";
            when "00" & x"3ed" => data <= x"05";
            when "00" & x"3ee" => data <= x"ba";
            when "00" & x"3ef" => data <= x"bd";
            when "00" & x"3f0" => data <= x"07";
            when "00" & x"3f1" => data <= x"01";
            when "00" & x"3f2" => data <= x"48";
            when "00" & x"3f3" => data <= x"88";
            when "00" & x"3f4" => data <= x"d0";
            when "00" & x"3f5" => data <= x"f8";
            when "00" & x"3f6" => data <= x"a0";
            when "00" & x"3f7" => data <= x"0a";
            when "00" & x"3f8" => data <= x"bd";
            when "00" & x"3f9" => data <= x"09";
            when "00" & x"3fa" => data <= x"01";
            when "00" & x"3fb" => data <= x"9d";
            when "00" & x"3fc" => data <= x"0b";
            when "00" & x"3fd" => data <= x"01";
            when "00" & x"3fe" => data <= x"ca";
            when "00" & x"3ff" => data <= x"88";
            when "00" & x"400" => data <= x"d0";
            when "00" & x"401" => data <= x"f6";
            when "00" & x"402" => data <= x"68";
            when "00" & x"403" => data <= x"68";
            when "00" & x"404" => data <= x"68";
            when "00" & x"405" => data <= x"a8";
            when "00" & x"406" => data <= x"68";
            when "00" & x"407" => data <= x"aa";
            when "00" & x"408" => data <= x"68";
            when "00" & x"409" => data <= x"60";
            when "00" & x"40a" => data <= x"ba";
            when "00" & x"40b" => data <= x"9d";
            when "00" & x"40c" => data <= x"03";
            when "00" & x"40d" => data <= x"01";
            when "00" & x"40e" => data <= x"4c";
            when "00" & x"40f" => data <= x"04";
            when "00" & x"410" => data <= x"84";
            when "00" & x"411" => data <= x"48";
            when "00" & x"412" => data <= x"8a";
            when "00" & x"413" => data <= x"48";
            when "00" & x"414" => data <= x"98";
            when "00" & x"415" => data <= x"48";
            when "00" & x"416" => data <= x"a9";
            when "00" & x"417" => data <= x"84";
            when "00" & x"418" => data <= x"48";
            when "00" & x"419" => data <= x"a9";
            when "00" & x"41a" => data <= x"09";
            when "00" & x"41b" => data <= x"48";
            when "00" & x"41c" => data <= x"d0";
            when "00" & x"41d" => data <= x"ce";
            when "00" & x"41e" => data <= x"20";
            when "00" & x"41f" => data <= x"b8";
            when "00" & x"420" => data <= x"86";
            when "00" & x"421" => data <= x"20";
            when "00" & x"422" => data <= x"3b";
            when "00" & x"423" => data <= x"af";
            when "00" & x"424" => data <= x"a0";
            when "00" & x"425" => data <= x"ff";
            when "00" & x"426" => data <= x"84";
            when "00" & x"427" => data <= x"a8";
            when "00" & x"428" => data <= x"c8";
            when "00" & x"429" => data <= x"84";
            when "00" & x"42a" => data <= x"aa";
            when "00" & x"42b" => data <= x"b9";
            when "00" & x"42c" => data <= x"00";
            when "00" & x"42d" => data <= x"0e";
            when "00" & x"42e" => data <= x"c0";
            when "00" & x"42f" => data <= x"08";
            when "00" & x"430" => data <= x"90";
            when "00" & x"431" => data <= x"03";
            when "00" & x"432" => data <= x"b9";
            when "00" & x"433" => data <= x"f8";
            when "00" & x"434" => data <= x"0e";
            when "00" & x"435" => data <= x"20";
            when "00" & x"436" => data <= x"9c";
            when "00" & x"437" => data <= x"80";
            when "00" & x"438" => data <= x"c8";
            when "00" & x"439" => data <= x"c0";
            when "00" & x"43a" => data <= x"0c";
            when "00" & x"43b" => data <= x"d0";
            when "00" & x"43c" => data <= x"ee";
            when "00" & x"43d" => data <= x"20";
            when "00" & x"43e" => data <= x"65";
            when "00" & x"43f" => data <= x"80";
            when "00" & x"440" => data <= x"20";
            when "00" & x"441" => data <= x"28";
            when "00" & x"442" => data <= x"ad";
            when "00" & x"443" => data <= x"04";
            when "00" & x"444" => data <= x"0f";
            when "00" & x"445" => data <= x"20";
            when "00" & x"446" => data <= x"c2";
            when "00" & x"447" => data <= x"80";
            when "00" & x"448" => data <= x"20";
            when "00" & x"449" => data <= x"65";
            when "00" & x"44a" => data <= x"80";
            when "00" & x"44b" => data <= x"29";
            when "00" & x"44c" => data <= x"0d";
            when "00" & x"44d" => data <= x"44";
            when "00" & x"44e" => data <= x"72";
            when "00" & x"44f" => data <= x"69";
            when "00" & x"450" => data <= x"76";
            when "00" & x"451" => data <= x"65";
            when "00" & x"452" => data <= x"20";
            when "00" & x"453" => data <= x"a5";
            when "00" & x"454" => data <= x"cf";
            when "00" & x"455" => data <= x"20";
            when "00" & x"456" => data <= x"ca";
            when "00" & x"457" => data <= x"80";
            when "00" & x"458" => data <= x"a0";
            when "00" & x"459" => data <= x"0d";
            when "00" & x"45a" => data <= x"20";
            when "00" & x"45b" => data <= x"f4";
            when "00" & x"45c" => data <= x"81";
            when "00" & x"45d" => data <= x"20";
            when "00" & x"45e" => data <= x"65";
            when "00" & x"45f" => data <= x"80";
            when "00" & x"460" => data <= x"4f";
            when "00" & x"461" => data <= x"70";
            when "00" & x"462" => data <= x"74";
            when "00" & x"463" => data <= x"69";
            when "00" & x"464" => data <= x"6f";
            when "00" & x"465" => data <= x"6e";
            when "00" & x"466" => data <= x"20";
            when "00" & x"467" => data <= x"ad";
            when "00" & x"468" => data <= x"06";
            when "00" & x"469" => data <= x"0f";
            when "00" & x"46a" => data <= x"20";
            when "00" & x"46b" => data <= x"05";
            when "00" & x"46c" => data <= x"82";
            when "00" & x"46d" => data <= x"20";
            when "00" & x"46e" => data <= x"ca";
            when "00" & x"46f" => data <= x"80";
            when "00" & x"470" => data <= x"20";
            when "00" & x"471" => data <= x"65";
            when "00" & x"472" => data <= x"80";
            when "00" & x"473" => data <= x"20";
            when "00" & x"474" => data <= x"28";
            when "00" & x"475" => data <= x"a0";
            when "00" & x"476" => data <= x"03";
            when "00" & x"477" => data <= x"0a";
            when "00" & x"478" => data <= x"0a";
            when "00" & x"479" => data <= x"aa";
            when "00" & x"47a" => data <= x"bd";
            when "00" & x"47b" => data <= x"6f";
            when "00" & x"47c" => data <= x"85";
            when "00" & x"47d" => data <= x"20";
            when "00" & x"47e" => data <= x"9c";
            when "00" & x"47f" => data <= x"80";
            when "00" & x"480" => data <= x"e8";
            when "00" & x"481" => data <= x"88";
            when "00" & x"482" => data <= x"10";
            when "00" & x"483" => data <= x"f6";
            when "00" & x"484" => data <= x"20";
            when "00" & x"485" => data <= x"65";
            when "00" & x"486" => data <= x"80";
            when "00" & x"487" => data <= x"29";
            when "00" & x"488" => data <= x"0d";
            when "00" & x"489" => data <= x"44";
            when "00" & x"48a" => data <= x"69";
            when "00" & x"48b" => data <= x"72";
            when "00" & x"48c" => data <= x"65";
            when "00" & x"48d" => data <= x"63";
            when "00" & x"48e" => data <= x"74";
            when "00" & x"48f" => data <= x"6f";
            when "00" & x"490" => data <= x"72";
            when "00" & x"491" => data <= x"79";
            when "00" & x"492" => data <= x"20";
            when "00" & x"493" => data <= x"3a";
            when "00" & x"494" => data <= x"ad";
            when "00" & x"495" => data <= x"cb";
            when "00" & x"496" => data <= x"10";
            when "00" & x"497" => data <= x"20";
            when "00" & x"498" => data <= x"ca";
            when "00" & x"499" => data <= x"80";
            when "00" & x"49a" => data <= x"20";
            when "00" & x"49b" => data <= x"9a";
            when "00" & x"49c" => data <= x"80";
            when "00" & x"49d" => data <= x"ad";
            when "00" & x"49e" => data <= x"ca";
            when "00" & x"49f" => data <= x"10";
            when "00" & x"4a0" => data <= x"20";
            when "00" & x"4a1" => data <= x"9c";
            when "00" & x"4a2" => data <= x"80";
            when "00" & x"4a3" => data <= x"a0";
            when "00" & x"4a4" => data <= x"06";
            when "00" & x"4a5" => data <= x"20";
            when "00" & x"4a6" => data <= x"f4";
            when "00" & x"4a7" => data <= x"81";
            when "00" & x"4a8" => data <= x"20";
            when "00" & x"4a9" => data <= x"65";
            when "00" & x"4aa" => data <= x"80";
            when "00" & x"4ab" => data <= x"4c";
            when "00" & x"4ac" => data <= x"69";
            when "00" & x"4ad" => data <= x"62";
            when "00" & x"4ae" => data <= x"72";
            when "00" & x"4af" => data <= x"61";
            when "00" & x"4b0" => data <= x"72";
            when "00" & x"4b1" => data <= x"79";
            when "00" & x"4b2" => data <= x"20";
            when "00" & x"4b3" => data <= x"3a";
            when "00" & x"4b4" => data <= x"ad";
            when "00" & x"4b5" => data <= x"cd";
            when "00" & x"4b6" => data <= x"10";
            when "00" & x"4b7" => data <= x"20";
            when "00" & x"4b8" => data <= x"ca";
            when "00" & x"4b9" => data <= x"80";
            when "00" & x"4ba" => data <= x"20";
            when "00" & x"4bb" => data <= x"9a";
            when "00" & x"4bc" => data <= x"80";
            when "00" & x"4bd" => data <= x"ad";
            when "00" & x"4be" => data <= x"cc";
            when "00" & x"4bf" => data <= x"10";
            when "00" & x"4c0" => data <= x"20";
            when "00" & x"4c1" => data <= x"9c";
            when "00" & x"4c2" => data <= x"80";
            when "00" & x"4c3" => data <= x"20";
            when "00" & x"4c4" => data <= x"9a";
            when "00" & x"4c5" => data <= x"9f";
            when "00" & x"4c6" => data <= x"a0";
            when "00" & x"4c7" => data <= x"00";
            when "00" & x"4c8" => data <= x"cc";
            when "00" & x"4c9" => data <= x"05";
            when "00" & x"4ca" => data <= x"0f";
            when "00" & x"4cb" => data <= x"b0";
            when "00" & x"4cc" => data <= x"17";
            when "00" & x"4cd" => data <= x"b9";
            when "00" & x"4ce" => data <= x"0f";
            when "00" & x"4cf" => data <= x"0e";
            when "00" & x"4d0" => data <= x"4d";
            when "00" & x"4d1" => data <= x"ca";
            when "00" & x"4d2" => data <= x"10";
            when "00" & x"4d3" => data <= x"29";
            when "00" & x"4d4" => data <= x"7f";
            when "00" & x"4d5" => data <= x"d0";
            when "00" & x"4d6" => data <= x"08";
            when "00" & x"4d7" => data <= x"b9";
            when "00" & x"4d8" => data <= x"0f";
            when "00" & x"4d9" => data <= x"0e";
            when "00" & x"4da" => data <= x"29";
            when "00" & x"4db" => data <= x"80";
            when "00" & x"4dc" => data <= x"99";
            when "00" & x"4dd" => data <= x"0f";
            when "00" & x"4de" => data <= x"0e";
            when "00" & x"4df" => data <= x"20";
            when "00" & x"4e0" => data <= x"10";
            when "00" & x"4e1" => data <= x"82";
            when "00" & x"4e2" => data <= x"90";
            when "00" & x"4e3" => data <= x"e4";
            when "00" & x"4e4" => data <= x"a0";
            when "00" & x"4e5" => data <= x"00";
            when "00" & x"4e6" => data <= x"20";
            when "00" & x"4e7" => data <= x"f6";
            when "00" & x"4e8" => data <= x"84";
            when "00" & x"4e9" => data <= x"90";
            when "00" & x"4ea" => data <= x"16";
            when "00" & x"4eb" => data <= x"a9";
            when "00" & x"4ec" => data <= x"ff";
            when "00" & x"4ed" => data <= x"8d";
            when "00" & x"4ee" => data <= x"82";
            when "00" & x"4ef" => data <= x"10";
            when "00" & x"4f0" => data <= x"4c";
            when "00" & x"4f1" => data <= x"9a";
            when "00" & x"4f2" => data <= x"9f";
            when "00" & x"4f3" => data <= x"20";
            when "00" & x"4f4" => data <= x"10";
            when "00" & x"4f5" => data <= x"82";
            when "00" & x"4f6" => data <= x"cc";
            when "00" & x"4f7" => data <= x"05";
            when "00" & x"4f8" => data <= x"0f";
            when "00" & x"4f9" => data <= x"b0";
            when "00" & x"4fa" => data <= x"05";
            when "00" & x"4fb" => data <= x"b9";
            when "00" & x"4fc" => data <= x"08";
            when "00" & x"4fd" => data <= x"0e";
            when "00" & x"4fe" => data <= x"30";
            when "00" & x"4ff" => data <= x"f3";
            when "00" & x"500" => data <= x"60";
            when "00" & x"501" => data <= x"84";
            when "00" & x"502" => data <= x"ab";
            when "00" & x"503" => data <= x"a2";
            when "00" & x"504" => data <= x"00";
            when "00" & x"505" => data <= x"b9";
            when "00" & x"506" => data <= x"08";
            when "00" & x"507" => data <= x"0e";
            when "00" & x"508" => data <= x"29";
            when "00" & x"509" => data <= x"7f";
            when "00" & x"50a" => data <= x"9d";
            when "00" & x"50b" => data <= x"60";
            when "00" & x"50c" => data <= x"10";
            when "00" & x"50d" => data <= x"c8";
            when "00" & x"50e" => data <= x"e8";
            when "00" & x"50f" => data <= x"e0";
            when "00" & x"510" => data <= x"08";
            when "00" & x"511" => data <= x"d0";
            when "00" & x"512" => data <= x"f2";
            when "00" & x"513" => data <= x"20";
            when "00" & x"514" => data <= x"f6";
            when "00" & x"515" => data <= x"84";
            when "00" & x"516" => data <= x"b0";
            when "00" & x"517" => data <= x"1f";
            when "00" & x"518" => data <= x"38";
            when "00" & x"519" => data <= x"a2";
            when "00" & x"51a" => data <= x"06";
            when "00" & x"51b" => data <= x"b9";
            when "00" & x"51c" => data <= x"0e";
            when "00" & x"51d" => data <= x"0e";
            when "00" & x"51e" => data <= x"fd";
            when "00" & x"51f" => data <= x"60";
            when "00" & x"520" => data <= x"10";
            when "00" & x"521" => data <= x"88";
            when "00" & x"522" => data <= x"ca";
            when "00" & x"523" => data <= x"10";
            when "00" & x"524" => data <= x"f6";
            when "00" & x"525" => data <= x"20";
            when "00" & x"526" => data <= x"11";
            when "00" & x"527" => data <= x"82";
            when "00" & x"528" => data <= x"b9";
            when "00" & x"529" => data <= x"0f";
            when "00" & x"52a" => data <= x"0e";
            when "00" & x"52b" => data <= x"29";
            when "00" & x"52c" => data <= x"7f";
            when "00" & x"52d" => data <= x"ed";
            when "00" & x"52e" => data <= x"67";
            when "00" & x"52f" => data <= x"10";
            when "00" & x"530" => data <= x"90";
            when "00" & x"531" => data <= x"cf";
            when "00" & x"532" => data <= x"20";
            when "00" & x"533" => data <= x"10";
            when "00" & x"534" => data <= x"82";
            when "00" & x"535" => data <= x"b0";
            when "00" & x"536" => data <= x"dc";
            when "00" & x"537" => data <= x"a4";
            when "00" & x"538" => data <= x"ab";
            when "00" & x"539" => data <= x"b9";
            when "00" & x"53a" => data <= x"08";
            when "00" & x"53b" => data <= x"0e";
            when "00" & x"53c" => data <= x"09";
            when "00" & x"53d" => data <= x"80";
            when "00" & x"53e" => data <= x"99";
            when "00" & x"53f" => data <= x"08";
            when "00" & x"540" => data <= x"0e";
            when "00" & x"541" => data <= x"ad";
            when "00" & x"542" => data <= x"67";
            when "00" & x"543" => data <= x"10";
            when "00" & x"544" => data <= x"c5";
            when "00" & x"545" => data <= x"aa";
            when "00" & x"546" => data <= x"f0";
            when "00" & x"547" => data <= x"10";
            when "00" & x"548" => data <= x"a6";
            when "00" & x"549" => data <= x"aa";
            when "00" & x"54a" => data <= x"85";
            when "00" & x"54b" => data <= x"aa";
            when "00" & x"54c" => data <= x"d0";
            when "00" & x"54d" => data <= x"0a";
            when "00" & x"54e" => data <= x"20";
            when "00" & x"54f" => data <= x"9a";
            when "00" & x"550" => data <= x"9f";
            when "00" & x"551" => data <= x"20";
            when "00" & x"552" => data <= x"9a";
            when "00" & x"553" => data <= x"9f";
            when "00" & x"554" => data <= x"a0";
            when "00" & x"555" => data <= x"ff";
            when "00" & x"556" => data <= x"d0";
            when "00" & x"557" => data <= x"09";
            when "00" & x"558" => data <= x"a4";
            when "00" & x"559" => data <= x"a8";
            when "00" & x"55a" => data <= x"d0";
            when "00" & x"55b" => data <= x"f5";
            when "00" & x"55c" => data <= x"a0";
            when "00" & x"55d" => data <= x"05";
            when "00" & x"55e" => data <= x"20";
            when "00" & x"55f" => data <= x"f4";
            when "00" & x"560" => data <= x"81";
            when "00" & x"561" => data <= x"c8";
            when "00" & x"562" => data <= x"84";
            when "00" & x"563" => data <= x"a8";
            when "00" & x"564" => data <= x"a4";
            when "00" & x"565" => data <= x"ab";
            when "00" & x"566" => data <= x"20";
            when "00" & x"567" => data <= x"cb";
            when "00" & x"568" => data <= x"9f";
            when "00" & x"569" => data <= x"20";
            when "00" & x"56a" => data <= x"c0";
            when "00" & x"56b" => data <= x"81";
            when "00" & x"56c" => data <= x"4c";
            when "00" & x"56d" => data <= x"e4";
            when "00" & x"56e" => data <= x"84";
            when "00" & x"56f" => data <= x"6f";
            when "00" & x"570" => data <= x"66";
            when "00" & x"571" => data <= x"66";
            when "00" & x"572" => data <= x"00";
            when "00" & x"573" => data <= x"4c";
            when "00" & x"574" => data <= x"4f";
            when "00" & x"575" => data <= x"41";
            when "00" & x"576" => data <= x"44";
            when "00" & x"577" => data <= x"52";
            when "00" & x"578" => data <= x"55";
            when "00" & x"579" => data <= x"4e";
            when "00" & x"57a" => data <= x"00";
            when "00" & x"57b" => data <= x"45";
            when "00" & x"57c" => data <= x"58";
            when "00" & x"57d" => data <= x"45";
            when "00" & x"57e" => data <= x"43";
            when "00" & x"57f" => data <= x"b9";
            when "00" & x"580" => data <= x"0e";
            when "00" & x"581" => data <= x"0f";
            when "00" & x"582" => data <= x"20";
            when "00" & x"583" => data <= x"fd";
            when "00" & x"584" => data <= x"81";
            when "00" & x"585" => data <= x"85";
            when "00" & x"586" => data <= x"c4";
            when "00" & x"587" => data <= x"18";
            when "00" & x"588" => data <= x"a9";
            when "00" & x"589" => data <= x"ff";
            when "00" & x"58a" => data <= x"79";
            when "00" & x"58b" => data <= x"0c";
            when "00" & x"58c" => data <= x"0f";
            when "00" & x"58d" => data <= x"b9";
            when "00" & x"58e" => data <= x"0f";
            when "00" & x"58f" => data <= x"0f";
            when "00" & x"590" => data <= x"79";
            when "00" & x"591" => data <= x"0d";
            when "00" & x"592" => data <= x"0f";
            when "00" & x"593" => data <= x"85";
            when "00" & x"594" => data <= x"c5";
            when "00" & x"595" => data <= x"b9";
            when "00" & x"596" => data <= x"0e";
            when "00" & x"597" => data <= x"0f";
            when "00" & x"598" => data <= x"29";
            when "00" & x"599" => data <= x"03";
            when "00" & x"59a" => data <= x"65";
            when "00" & x"59b" => data <= x"c4";
            when "00" & x"59c" => data <= x"85";
            when "00" & x"59d" => data <= x"c4";
            when "00" & x"59e" => data <= x"38";
            when "00" & x"59f" => data <= x"b9";
            when "00" & x"5a0" => data <= x"07";
            when "00" & x"5a1" => data <= x"0f";
            when "00" & x"5a2" => data <= x"e5";
            when "00" & x"5a3" => data <= x"c5";
            when "00" & x"5a4" => data <= x"48";
            when "00" & x"5a5" => data <= x"b9";
            when "00" & x"5a6" => data <= x"06";
            when "00" & x"5a7" => data <= x"0f";
            when "00" & x"5a8" => data <= x"29";
            when "00" & x"5a9" => data <= x"03";
            when "00" & x"5aa" => data <= x"e5";
            when "00" & x"5ab" => data <= x"c4";
            when "00" & x"5ac" => data <= x"aa";
            when "00" & x"5ad" => data <= x"a9";
            when "00" & x"5ae" => data <= x"00";
            when "00" & x"5af" => data <= x"c5";
            when "00" & x"5b0" => data <= x"c2";
            when "00" & x"5b1" => data <= x"68";
            when "00" & x"5b2" => data <= x"e5";
            when "00" & x"5b3" => data <= x"c3";
            when "00" & x"5b4" => data <= x"8a";
            when "00" & x"5b5" => data <= x"e5";
            when "00" & x"5b6" => data <= x"c6";
            when "00" & x"5b7" => data <= x"60";
            when "00" & x"5b8" => data <= x"41";
            when "00" & x"5b9" => data <= x"43";
            when "00" & x"5ba" => data <= x"43";
            when "00" & x"5bb" => data <= x"45";
            when "00" & x"5bc" => data <= x"53";
            when "00" & x"5bd" => data <= x"53";
            when "00" & x"5be" => data <= x"88";
            when "00" & x"5bf" => data <= x"d1";
            when "00" & x"5c0" => data <= x"32";
            when "00" & x"5c1" => data <= x"42";
            when "00" & x"5c2" => data <= x"41";
            when "00" & x"5c3" => data <= x"43";
            when "00" & x"5c4" => data <= x"4b";
            when "00" & x"5c5" => data <= x"55";
            when "00" & x"5c6" => data <= x"50";
            when "00" & x"5c7" => data <= x"9c";
            when "00" & x"5c8" => data <= x"ba";
            when "00" & x"5c9" => data <= x"54";
            when "00" & x"5ca" => data <= x"43";
            when "00" & x"5cb" => data <= x"4f";
            when "00" & x"5cc" => data <= x"4d";
            when "00" & x"5cd" => data <= x"50";
            when "00" & x"5ce" => data <= x"41";
            when "00" & x"5cf" => data <= x"43";
            when "00" & x"5d0" => data <= x"54";
            when "00" & x"5d1" => data <= x"9a";
            when "00" & x"5d2" => data <= x"bf";
            when "00" & x"5d3" => data <= x"0a";
            when "00" & x"5d4" => data <= x"43";
            when "00" & x"5d5" => data <= x"4f";
            when "00" & x"5d6" => data <= x"50";
            when "00" & x"5d7" => data <= x"59";
            when "00" & x"5d8" => data <= x"9d";
            when "00" & x"5d9" => data <= x"26";
            when "00" & x"5da" => data <= x"64";
            when "00" & x"5db" => data <= x"44";
            when "00" & x"5dc" => data <= x"45";
            when "00" & x"5dd" => data <= x"4c";
            when "00" & x"5de" => data <= x"45";
            when "00" & x"5df" => data <= x"54";
            when "00" & x"5e0" => data <= x"45";
            when "00" & x"5e1" => data <= x"86";
            when "00" & x"5e2" => data <= x"fd";
            when "00" & x"5e3" => data <= x"01";
            when "00" & x"5e4" => data <= x"44";
            when "00" & x"5e5" => data <= x"45";
            when "00" & x"5e6" => data <= x"53";
            when "00" & x"5e7" => data <= x"54";
            when "00" & x"5e8" => data <= x"52";
            when "00" & x"5e9" => data <= x"4f";
            when "00" & x"5ea" => data <= x"59";
            when "00" & x"5eb" => data <= x"87";
            when "00" & x"5ec" => data <= x"0f";
            when "00" & x"5ed" => data <= x"02";
            when "00" & x"5ee" => data <= x"44";
            when "00" & x"5ef" => data <= x"49";
            when "00" & x"5f0" => data <= x"52";
            when "00" & x"5f1" => data <= x"88";
            when "00" & x"5f2" => data <= x"4d";
            when "00" & x"5f3" => data <= x"09";
            when "00" & x"5f4" => data <= x"44";
            when "00" & x"5f5" => data <= x"52";
            when "00" & x"5f6" => data <= x"49";
            when "00" & x"5f7" => data <= x"56";
            when "00" & x"5f8" => data <= x"45";
            when "00" & x"5f9" => data <= x"87";
            when "00" & x"5fa" => data <= x"74";
            when "00" & x"5fb" => data <= x"0a";
            when "00" & x"5fc" => data <= x"45";
            when "00" & x"5fd" => data <= x"4e";
            when "00" & x"5fe" => data <= x"41";
            when "00" & x"5ff" => data <= x"42";
            when "00" & x"600" => data <= x"4c";
            when "00" & x"601" => data <= x"45";
            when "00" & x"602" => data <= x"8a";
            when "00" & x"603" => data <= x"38";
            when "00" & x"604" => data <= x"00";
            when "00" & x"605" => data <= x"49";
            when "00" & x"606" => data <= x"4e";
            when "00" & x"607" => data <= x"46";
            when "00" & x"608" => data <= x"4f";
            when "00" & x"609" => data <= x"82";
            when "00" & x"60a" => data <= x"83";
            when "00" & x"60b" => data <= x"02";
            when "00" & x"60c" => data <= x"4c";
            when "00" & x"60d" => data <= x"49";
            when "00" & x"60e" => data <= x"42";
            when "00" & x"60f" => data <= x"88";
            when "00" & x"610" => data <= x"51";
            when "00" & x"611" => data <= x"09";
            when "00" & x"612" => data <= x"52";
            when "00" & x"613" => data <= x"45";
            when "00" & x"614" => data <= x"4e";
            when "00" & x"615" => data <= x"41";
            when "00" & x"616" => data <= x"4d";
            when "00" & x"617" => data <= x"45";
            when "00" & x"618" => data <= x"8a";
            when "00" & x"619" => data <= x"6c";
            when "00" & x"61a" => data <= x"87";
            when "00" & x"61b" => data <= x"54";
            when "00" & x"61c" => data <= x"49";
            when "00" & x"61d" => data <= x"54";
            when "00" & x"61e" => data <= x"4c";
            when "00" & x"61f" => data <= x"45";
            when "00" & x"620" => data <= x"88";
            when "00" & x"621" => data <= x"a2";
            when "00" & x"622" => data <= x"0b";
            when "00" & x"623" => data <= x"57";
            when "00" & x"624" => data <= x"49";
            when "00" & x"625" => data <= x"50";
            when "00" & x"626" => data <= x"45";
            when "00" & x"627" => data <= x"86";
            when "00" & x"628" => data <= x"c2";
            when "00" & x"629" => data <= x"02";
            when "00" & x"62a" => data <= x"b4";
            when "00" & x"62b" => data <= x"6b";
            when "00" & x"62c" => data <= x"00";
            when "00" & x"62d" => data <= x"42";
            when "00" & x"62e" => data <= x"55";
            when "00" & x"62f" => data <= x"49";
            when "00" & x"630" => data <= x"4c";
            when "00" & x"631" => data <= x"44";
            when "00" & x"632" => data <= x"9f";
            when "00" & x"633" => data <= x"47";
            when "00" & x"634" => data <= x"01";
            when "00" & x"635" => data <= x"43";
            when "00" & x"636" => data <= x"41";
            when "00" & x"637" => data <= x"52";
            when "00" & x"638" => data <= x"44";
            when "00" & x"639" => data <= x"93";
            when "00" & x"63a" => data <= x"37";
            when "00" & x"63b" => data <= x"00";
            when "00" & x"63c" => data <= x"44";
            when "00" & x"63d" => data <= x"55";
            when "00" & x"63e" => data <= x"4d";
            when "00" & x"63f" => data <= x"50";
            when "00" & x"640" => data <= x"9e";
            when "00" & x"641" => data <= x"cf";
            when "00" & x"642" => data <= x"01";
            when "00" & x"643" => data <= x"4c";
            when "00" & x"644" => data <= x"49";
            when "00" & x"645" => data <= x"53";
            when "00" & x"646" => data <= x"54";
            when "00" & x"647" => data <= x"9e";
            when "00" & x"648" => data <= x"8d";
            when "00" & x"649" => data <= x"01";
            when "00" & x"64a" => data <= x"54";
            when "00" & x"64b" => data <= x"59";
            when "00" & x"64c" => data <= x"50";
            when "00" & x"64d" => data <= x"45";
            when "00" & x"64e" => data <= x"9e";
            when "00" & x"64f" => data <= x"86";
            when "00" & x"650" => data <= x"01";
            when "00" & x"651" => data <= x"44";
            when "00" & x"652" => data <= x"4d";
            when "00" & x"653" => data <= x"4d";
            when "00" & x"654" => data <= x"43";
            when "00" & x"655" => data <= x"93";
            when "00" & x"656" => data <= x"37";
            when "00" & x"657" => data <= x"00";
            when "00" & x"658" => data <= x"85";
            when "00" & x"659" => data <= x"b6";
            when "00" & x"65a" => data <= x"00";
            when "00" & x"65b" => data <= x"44";
            when "00" & x"65c" => data <= x"46";
            when "00" & x"65d" => data <= x"53";
            when "00" & x"65e" => data <= x"99";
            when "00" & x"65f" => data <= x"c5";
            when "00" & x"660" => data <= x"00";
            when "00" & x"661" => data <= x"55";
            when "00" & x"662" => data <= x"54";
            when "00" & x"663" => data <= x"49";
            when "00" & x"664" => data <= x"4c";
            when "00" & x"665" => data <= x"53";
            when "00" & x"666" => data <= x"99";
            when "00" & x"667" => data <= x"ed";
            when "00" & x"668" => data <= x"00";
            when "00" & x"669" => data <= x"99";
            when "00" & x"66a" => data <= x"f4";
            when "00" & x"66b" => data <= x"00";
            when "00" & x"66c" => data <= x"20";
            when "00" & x"66d" => data <= x"b8";
            when "00" & x"66e" => data <= x"86";
            when "00" & x"66f" => data <= x"a2";
            when "00" & x"670" => data <= x"fd";
            when "00" & x"671" => data <= x"8a";
            when "00" & x"672" => data <= x"ba";
            when "00" & x"673" => data <= x"86";
            when "00" & x"674" => data <= x"b6";
            when "00" & x"675" => data <= x"aa";
            when "00" & x"676" => data <= x"98";
            when "00" & x"677" => data <= x"48";
            when "00" & x"678" => data <= x"e8";
            when "00" & x"679" => data <= x"e8";
            when "00" & x"67a" => data <= x"68";
            when "00" & x"67b" => data <= x"48";
            when "00" & x"67c" => data <= x"a8";
            when "00" & x"67d" => data <= x"20";
            when "00" & x"67e" => data <= x"bf";
            when "00" & x"67f" => data <= x"86";
            when "00" & x"680" => data <= x"e8";
            when "00" & x"681" => data <= x"bd";
            when "00" & x"682" => data <= x"b8";
            when "00" & x"683" => data <= x"85";
            when "00" & x"684" => data <= x"30";
            when "00" & x"685" => data <= x"28";
            when "00" & x"686" => data <= x"ca";
            when "00" & x"687" => data <= x"88";
            when "00" & x"688" => data <= x"86";
            when "00" & x"689" => data <= x"b8";
            when "00" & x"68a" => data <= x"e8";
            when "00" & x"68b" => data <= x"c8";
            when "00" & x"68c" => data <= x"bd";
            when "00" & x"68d" => data <= x"b8";
            when "00" & x"68e" => data <= x"85";
            when "00" & x"68f" => data <= x"30";
            when "00" & x"690" => data <= x"16";
            when "00" & x"691" => data <= x"51";
            when "00" & x"692" => data <= x"f2";
            when "00" & x"693" => data <= x"29";
            when "00" & x"694" => data <= x"5f";
            when "00" & x"695" => data <= x"f0";
            when "00" & x"696" => data <= x"f3";
            when "00" & x"697" => data <= x"ca";
            when "00" & x"698" => data <= x"e8";
            when "00" & x"699" => data <= x"bd";
            when "00" & x"69a" => data <= x"b8";
            when "00" & x"69b" => data <= x"85";
            when "00" & x"69c" => data <= x"10";
            when "00" & x"69d" => data <= x"fa";
            when "00" & x"69e" => data <= x"b1";
            when "00" & x"69f" => data <= x"f2";
            when "00" & x"6a0" => data <= x"c9";
            when "00" & x"6a1" => data <= x"2e";
            when "00" & x"6a2" => data <= x"d0";
            when "00" & x"6a3" => data <= x"d4";
            when "00" & x"6a4" => data <= x"c8";
            when "00" & x"6a5" => data <= x"b0";
            when "00" & x"6a6" => data <= x"07";
            when "00" & x"6a7" => data <= x"b1";
            when "00" & x"6a8" => data <= x"f2";
            when "00" & x"6a9" => data <= x"20";
            when "00" & x"6aa" => data <= x"ee";
            when "00" & x"6ab" => data <= x"82";
            when "00" & x"6ac" => data <= x"90";
            when "00" & x"6ad" => data <= x"ca";
            when "00" & x"6ae" => data <= x"68";
            when "00" & x"6af" => data <= x"bd";
            when "00" & x"6b0" => data <= x"b8";
            when "00" & x"6b1" => data <= x"85";
            when "00" & x"6b2" => data <= x"48";
            when "00" & x"6b3" => data <= x"bd";
            when "00" & x"6b4" => data <= x"b9";
            when "00" & x"6b5" => data <= x"85";
            when "00" & x"6b6" => data <= x"48";
            when "00" & x"6b7" => data <= x"60";
            when "00" & x"6b8" => data <= x"86";
            when "00" & x"6b9" => data <= x"f2";
            when "00" & x"6ba" => data <= x"84";
            when "00" & x"6bb" => data <= x"f3";
            when "00" & x"6bc" => data <= x"a0";
            when "00" & x"6bd" => data <= x"00";
            when "00" & x"6be" => data <= x"60";
            when "00" & x"6bf" => data <= x"18";
            when "00" & x"6c0" => data <= x"4c";
            when "00" & x"6c1" => data <= x"c2";
            when "00" & x"6c2" => data <= x"ff";
            when "00" & x"6c3" => data <= x"20";
            when "00" & x"6c4" => data <= x"5e";
            when "00" & x"6c5" => data <= x"82";
            when "00" & x"6c6" => data <= x"20";
            when "00" & x"6c7" => data <= x"01";
            when "00" & x"6c8" => data <= x"9a";
            when "00" & x"6c9" => data <= x"20";
            when "00" & x"6ca" => data <= x"68";
            when "00" & x"6cb" => data <= x"82";
            when "00" & x"6cc" => data <= x"b9";
            when "00" & x"6cd" => data <= x"0f";
            when "00" & x"6ce" => data <= x"0e";
            when "00" & x"6cf" => data <= x"30";
            when "00" & x"6d0" => data <= x"12";
            when "00" & x"6d1" => data <= x"20";
            when "00" & x"6d2" => data <= x"c0";
            when "00" & x"6d3" => data <= x"81";
            when "00" & x"6d4" => data <= x"20";
            when "00" & x"6d5" => data <= x"65";
            when "00" & x"6d6" => data <= x"80";
            when "00" & x"6d7" => data <= x"20";
            when "00" & x"6d8" => data <= x"3a";
            when "00" & x"6d9" => data <= x"20";
            when "00" & x"6da" => data <= x"ea";
            when "00" & x"6db" => data <= x"20";
            when "00" & x"6dc" => data <= x"9e";
            when "00" & x"6dd" => data <= x"9c";
            when "00" & x"6de" => data <= x"f0";
            when "00" & x"6df" => data <= x"09";
            when "00" & x"6e0" => data <= x"20";
            when "00" & x"6e1" => data <= x"9a";
            when "00" & x"6e2" => data <= x"9f";
            when "00" & x"6e3" => data <= x"20";
            when "00" & x"6e4" => data <= x"9d";
            when "00" & x"6e5" => data <= x"82";
            when "00" & x"6e6" => data <= x"b0";
            when "00" & x"6e7" => data <= x"e4";
            when "00" & x"6e8" => data <= x"60";
            when "00" & x"6e9" => data <= x"20";
            when "00" & x"6ea" => data <= x"a1";
            when "00" & x"6eb" => data <= x"81";
            when "00" & x"6ec" => data <= x"20";
            when "00" & x"6ed" => data <= x"d1";
            when "00" & x"6ee" => data <= x"82";
            when "00" & x"6ef" => data <= x"20";
            when "00" & x"6f0" => data <= x"b4";
            when "00" & x"6f1" => data <= x"8a";
            when "00" & x"6f2" => data <= x"ac";
            when "00" & x"6f3" => data <= x"ce";
            when "00" & x"6f4" => data <= x"10";
            when "00" & x"6f5" => data <= x"20";
            when "00" & x"6f6" => data <= x"19";
            when "00" & x"6f7" => data <= x"82";
            when "00" & x"6f8" => data <= x"8c";
            when "00" & x"6f9" => data <= x"ce";
            when "00" & x"6fa" => data <= x"10";
            when "00" & x"6fb" => data <= x"4c";
            when "00" & x"6fc" => data <= x"e0";
            when "00" & x"6fd" => data <= x"86";
            when "00" & x"6fe" => data <= x"20";
            when "00" & x"6ff" => data <= x"62";
            when "00" & x"700" => data <= x"82";
            when "00" & x"701" => data <= x"20";
            when "00" & x"702" => data <= x"01";
            when "00" & x"703" => data <= x"9a";
            when "00" & x"704" => data <= x"20";
            when "00" & x"705" => data <= x"68";
            when "00" & x"706" => data <= x"82";
            when "00" & x"707" => data <= x"20";
            when "00" & x"708" => data <= x"fc";
            when "00" & x"709" => data <= x"82";
            when "00" & x"70a" => data <= x"20";
            when "00" & x"70b" => data <= x"d1";
            when "00" & x"70c" => data <= x"82";
            when "00" & x"70d" => data <= x"4c";
            when "00" & x"70e" => data <= x"b4";
            when "00" & x"70f" => data <= x"8a";
            when "00" & x"710" => data <= x"20";
            when "00" & x"711" => data <= x"bd";
            when "00" & x"712" => data <= x"9b";
            when "00" & x"713" => data <= x"20";
            when "00" & x"714" => data <= x"5e";
            when "00" & x"715" => data <= x"82";
            when "00" & x"716" => data <= x"20";
            when "00" & x"717" => data <= x"01";
            when "00" & x"718" => data <= x"9a";
            when "00" & x"719" => data <= x"20";
            when "00" & x"71a" => data <= x"68";
            when "00" & x"71b" => data <= x"82";
            when "00" & x"71c" => data <= x"b9";
            when "00" & x"71d" => data <= x"0f";
            when "00" & x"71e" => data <= x"0e";
            when "00" & x"71f" => data <= x"30";
            when "00" & x"720" => data <= x"06";
            when "00" & x"721" => data <= x"20";
            when "00" & x"722" => data <= x"c0";
            when "00" & x"723" => data <= x"81";
            when "00" & x"724" => data <= x"20";
            when "00" & x"725" => data <= x"9a";
            when "00" & x"726" => data <= x"9f";
            when "00" & x"727" => data <= x"20";
            when "00" & x"728" => data <= x"9d";
            when "00" & x"729" => data <= x"82";
            when "00" & x"72a" => data <= x"b0";
            when "00" & x"72b" => data <= x"f0";
            when "00" & x"72c" => data <= x"20";
            when "00" & x"72d" => data <= x"65";
            when "00" & x"72e" => data <= x"80";
            when "00" & x"72f" => data <= x"0d";
            when "00" & x"730" => data <= x"44";
            when "00" & x"731" => data <= x"65";
            when "00" & x"732" => data <= x"6c";
            when "00" & x"733" => data <= x"65";
            when "00" & x"734" => data <= x"74";
            when "00" & x"735" => data <= x"65";
            when "00" & x"736" => data <= x"20";
            when "00" & x"737" => data <= x"28";
            when "00" & x"738" => data <= x"59";
            when "00" & x"739" => data <= x"2f";
            when "00" & x"73a" => data <= x"4e";
            when "00" & x"73b" => data <= x"29";
            when "00" & x"73c" => data <= x"20";
            when "00" & x"73d" => data <= x"3f";
            when "00" & x"73e" => data <= x"20";
            when "00" & x"73f" => data <= x"ea";
            when "00" & x"740" => data <= x"20";
            when "00" & x"741" => data <= x"9e";
            when "00" & x"742" => data <= x"9c";
            when "00" & x"743" => data <= x"f0";
            when "00" & x"744" => data <= x"03";
            when "00" & x"745" => data <= x"4c";
            when "00" & x"746" => data <= x"9a";
            when "00" & x"747" => data <= x"9f";
            when "00" & x"748" => data <= x"20";
            when "00" & x"749" => data <= x"a1";
            when "00" & x"74a" => data <= x"81";
            when "00" & x"74b" => data <= x"20";
            when "00" & x"74c" => data <= x"96";
            when "00" & x"74d" => data <= x"82";
            when "00" & x"74e" => data <= x"b9";
            when "00" & x"74f" => data <= x"0f";
            when "00" & x"750" => data <= x"0e";
            when "00" & x"751" => data <= x"30";
            when "00" & x"752" => data <= x"0c";
            when "00" & x"753" => data <= x"20";
            when "00" & x"754" => data <= x"d1";
            when "00" & x"755" => data <= x"82";
            when "00" & x"756" => data <= x"ac";
            when "00" & x"757" => data <= x"ce";
            when "00" & x"758" => data <= x"10";
            when "00" & x"759" => data <= x"20";
            when "00" & x"75a" => data <= x"19";
            when "00" & x"75b" => data <= x"82";
            when "00" & x"75c" => data <= x"8c";
            when "00" & x"75d" => data <= x"ce";
            when "00" & x"75e" => data <= x"10";
            when "00" & x"75f" => data <= x"20";
            when "00" & x"760" => data <= x"9d";
            when "00" & x"761" => data <= x"82";
            when "00" & x"762" => data <= x"b0";
            when "00" & x"763" => data <= x"ea";
            when "00" & x"764" => data <= x"20";
            when "00" & x"765" => data <= x"b4";
            when "00" & x"766" => data <= x"8a";
            when "00" & x"767" => data <= x"20";
            when "00" & x"768" => data <= x"65";
            when "00" & x"769" => data <= x"80";
            when "00" & x"76a" => data <= x"0d";
            when "00" & x"76b" => data <= x"44";
            when "00" & x"76c" => data <= x"65";
            when "00" & x"76d" => data <= x"6c";
            when "00" & x"76e" => data <= x"65";
            when "00" & x"76f" => data <= x"74";
            when "00" & x"770" => data <= x"65";
            when "00" & x"771" => data <= x"64";
            when "00" & x"772" => data <= x"0d";
            when "00" & x"773" => data <= x"ea";
            when "00" & x"774" => data <= x"60";
            when "00" & x"775" => data <= x"20";
            when "00" & x"776" => data <= x"01";
            when "00" & x"777" => data <= x"9a";
            when "00" & x"778" => data <= x"20";
            when "00" & x"779" => data <= x"5d";
            when "00" & x"77a" => data <= x"83";
            when "00" & x"77b" => data <= x"8d";
            when "00" & x"77c" => data <= x"cb";
            when "00" & x"77d" => data <= x"10";
            when "00" & x"77e" => data <= x"ea";
            when "00" & x"77f" => data <= x"ea";
            when "00" & x"780" => data <= x"ea";
            when "00" & x"781" => data <= x"29";
            when "00" & x"782" => data <= x"03";
            when "00" & x"783" => data <= x"85";
            when "00" & x"784" => data <= x"cf";
            when "00" & x"785" => data <= x"60";
            when "00" & x"786" => data <= x"20";
            when "00" & x"787" => data <= x"61";
            when "00" & x"788" => data <= x"89";
            when "00" & x"789" => data <= x"20";
            when "00" & x"78a" => data <= x"6e";
            when "00" & x"78b" => data <= x"98";
            when "00" & x"78c" => data <= x"20";
            when "00" & x"78d" => data <= x"7e";
            when "00" & x"78e" => data <= x"83";
            when "00" & x"78f" => data <= x"4c";
            when "00" & x"790" => data <= x"99";
            when "00" & x"791" => data <= x"af";
            when "00" & x"792" => data <= x"ea";
            when "00" & x"793" => data <= x"ea";
            when "00" & x"794" => data <= x"20";
            when "00" & x"795" => data <= x"6e";
            when "00" & x"796" => data <= x"82";
            when "00" & x"797" => data <= x"20";
            when "00" & x"798" => data <= x"6e";
            when "00" & x"799" => data <= x"98";
            when "00" & x"79a" => data <= x"20";
            when "00" & x"79b" => data <= x"7e";
            when "00" & x"79c" => data <= x"83";
            when "00" & x"79d" => data <= x"84";
            when "00" & x"79e" => data <= x"bc";
            when "00" & x"79f" => data <= x"a2";
            when "00" & x"7a0" => data <= x"00";
            when "00" & x"7a1" => data <= x"a5";
            when "00" & x"7a2" => data <= x"c0";
            when "00" & x"7a3" => data <= x"d0";
            when "00" & x"7a4" => data <= x"06";
            when "00" & x"7a5" => data <= x"c8";
            when "00" & x"7a6" => data <= x"c8";
            when "00" & x"7a7" => data <= x"a2";
            when "00" & x"7a8" => data <= x"02";
            when "00" & x"7a9" => data <= x"d0";
            when "00" & x"7aa" => data <= x"08";
            when "00" & x"7ab" => data <= x"b9";
            when "00" & x"7ac" => data <= x"0e";
            when "00" & x"7ad" => data <= x"0f";
            when "00" & x"7ae" => data <= x"85";
            when "00" & x"7af" => data <= x"c4";
            when "00" & x"7b0" => data <= x"20";
            when "00" & x"7b1" => data <= x"3f";
            when "00" & x"7b2" => data <= x"8a";
            when "00" & x"7b3" => data <= x"b9";
            when "00" & x"7b4" => data <= x"08";
            when "00" & x"7b5" => data <= x"0f";
            when "00" & x"7b6" => data <= x"95";
            when "00" & x"7b7" => data <= x"be";
            when "00" & x"7b8" => data <= x"c8";
            when "00" & x"7b9" => data <= x"e8";
            when "00" & x"7ba" => data <= x"e0";
            when "00" & x"7bb" => data <= x"08";
            when "00" & x"7bc" => data <= x"d0";
            when "00" & x"7bd" => data <= x"f5";
            when "00" & x"7be" => data <= x"20";
            when "00" & x"7bf" => data <= x"56";
            when "00" & x"7c0" => data <= x"8a";
            when "00" & x"7c1" => data <= x"a4";
            when "00" & x"7c2" => data <= x"bc";
            when "00" & x"7c3" => data <= x"20";
            when "00" & x"7c4" => data <= x"fc";
            when "00" & x"7c5" => data <= x"82";
            when "00" & x"7c6" => data <= x"4c";
            when "00" & x"7c7" => data <= x"8a";
            when "00" & x"7c8" => data <= x"af";
            when "00" & x"7c9" => data <= x"00";
            when "00" & x"7ca" => data <= x"00";
            when "00" & x"7cb" => data <= x"00";
            when "00" & x"7cc" => data <= x"00";
            when "00" & x"7cd" => data <= x"00";
            when "00" & x"7ce" => data <= x"00";
            when "00" & x"7cf" => data <= x"00";
            when "00" & x"7d0" => data <= x"00";
            when "00" & x"7d1" => data <= x"00";
            when "00" & x"7d2" => data <= x"00";
            when "00" & x"7d3" => data <= x"00";
            when "00" & x"7d4" => data <= x"20";
            when "00" & x"7d5" => data <= x"b8";
            when "00" & x"7d6" => data <= x"86";
            when "00" & x"7d7" => data <= x"20";
            when "00" & x"7d8" => data <= x"41";
            when "00" & x"7d9" => data <= x"88";
            when "00" & x"7da" => data <= x"8c";
            when "00" & x"7db" => data <= x"db";
            when "00" & x"7dc" => data <= x"10";
            when "00" & x"7dd" => data <= x"20";
            when "00" & x"7de" => data <= x"06";
            when "00" & x"7df" => data <= x"81";
            when "00" & x"7e0" => data <= x"8c";
            when "00" & x"7e1" => data <= x"da";
            when "00" & x"7e2" => data <= x"10";
            when "00" & x"7e3" => data <= x"20";
            when "00" & x"7e4" => data <= x"96";
            when "00" & x"7e5" => data <= x"82";
            when "00" & x"7e6" => data <= x"b0";
            when "00" & x"7e7" => data <= x"22";
            when "00" & x"7e8" => data <= x"ac";
            when "00" & x"7e9" => data <= x"db";
            when "00" & x"7ea" => data <= x"10";
            when "00" & x"7eb" => data <= x"ad";
            when "00" & x"7ec" => data <= x"cc";
            when "00" & x"7ed" => data <= x"10";
            when "00" & x"7ee" => data <= x"85";
            when "00" & x"7ef" => data <= x"ce";
            when "00" & x"7f0" => data <= x"ad";
            when "00" & x"7f1" => data <= x"cd";
            when "00" & x"7f2" => data <= x"10";
            when "00" & x"7f3" => data <= x"20";
            when "00" & x"7f4" => data <= x"7e";
            when "00" & x"7f5" => data <= x"87";
            when "00" & x"7f6" => data <= x"20";
            when "00" & x"7f7" => data <= x"09";
            when "00" & x"7f8" => data <= x"81";
            when "00" & x"7f9" => data <= x"20";
            when "00" & x"7fa" => data <= x"96";
            when "00" & x"7fb" => data <= x"82";
            when "00" & x"7fc" => data <= x"b0";
            when "00" & x"7fd" => data <= x"0c";
            when "00" & x"7fe" => data <= x"20";
            when "00" & x"7ff" => data <= x"22";
            when "00" & x"800" => data <= x"80";
            when "00" & x"801" => data <= x"fe";
            when "00" & x"802" => data <= x"63";
            when "00" & x"803" => data <= x"6f";
            when "00" & x"804" => data <= x"6d";
            when "00" & x"805" => data <= x"6d";
            when "00" & x"806" => data <= x"61";
            when "00" & x"807" => data <= x"6e";
            when "00" & x"808" => data <= x"64";
            when "00" & x"809" => data <= x"00";
            when "00" & x"80a" => data <= x"20";
            when "00" & x"80b" => data <= x"9d";
            when "00" & x"80c" => data <= x"87";
            when "00" & x"80d" => data <= x"18";
            when "00" & x"80e" => data <= x"ad";
            when "00" & x"80f" => data <= x"da";
            when "00" & x"810" => data <= x"10";
            when "00" & x"811" => data <= x"a8";
            when "00" & x"812" => data <= x"65";
            when "00" & x"813" => data <= x"f2";
            when "00" & x"814" => data <= x"8d";
            when "00" & x"815" => data <= x"da";
            when "00" & x"816" => data <= x"10";
            when "00" & x"817" => data <= x"a5";
            when "00" & x"818" => data <= x"f3";
            when "00" & x"819" => data <= x"69";
            when "00" & x"81a" => data <= x"00";
            when "00" & x"81b" => data <= x"8d";
            when "00" & x"81c" => data <= x"db";
            when "00" & x"81d" => data <= x"10";
            when "00" & x"81e" => data <= x"ad";
            when "00" & x"81f" => data <= x"76";
            when "00" & x"820" => data <= x"10";
            when "00" & x"821" => data <= x"2d";
            when "00" & x"822" => data <= x"77";
            when "00" & x"823" => data <= x"10";
            when "00" & x"824" => data <= x"0d";
            when "00" & x"825" => data <= x"d7";
            when "00" & x"826" => data <= x"10";
            when "00" & x"827" => data <= x"c9";
            when "00" & x"828" => data <= x"ff";
            when "00" & x"829" => data <= x"f0";
            when "00" & x"82a" => data <= x"13";
            when "00" & x"82b" => data <= x"a5";
            when "00" & x"82c" => data <= x"c0";
            when "00" & x"82d" => data <= x"8d";
            when "00" & x"82e" => data <= x"74";
            when "00" & x"82f" => data <= x"10";
            when "00" & x"830" => data <= x"a5";
            when "00" & x"831" => data <= x"c1";
            when "00" & x"832" => data <= x"8d";
            when "00" & x"833" => data <= x"75";
            when "00" & x"834" => data <= x"10";
            when "00" & x"835" => data <= x"a2";
            when "00" & x"836" => data <= x"74";
            when "00" & x"837" => data <= x"a0";
            when "00" & x"838" => data <= x"10";
            when "00" & x"839" => data <= x"a9";
            when "00" & x"83a" => data <= x"04";
            when "00" & x"83b" => data <= x"4c";
            when "00" & x"83c" => data <= x"06";
            when "00" & x"83d" => data <= x"04";
            when "00" & x"83e" => data <= x"6c";
            when "00" & x"83f" => data <= x"c0";
            when "00" & x"840" => data <= x"00";
            when "00" & x"841" => data <= x"a9";
            when "00" & x"842" => data <= x"ff";
            when "00" & x"843" => data <= x"85";
            when "00" & x"844" => data <= x"c0";
            when "00" & x"845" => data <= x"a5";
            when "00" & x"846" => data <= x"f2";
            when "00" & x"847" => data <= x"85";
            when "00" & x"848" => data <= x"bc";
            when "00" & x"849" => data <= x"a5";
            when "00" & x"84a" => data <= x"f3";
            when "00" & x"84b" => data <= x"85";
            when "00" & x"84c" => data <= x"bd";
            when "00" & x"84d" => data <= x"60";
            when "00" & x"84e" => data <= x"a2";
            when "00" & x"84f" => data <= x"00";
            when "00" & x"850" => data <= x"f0";
            when "00" & x"851" => data <= x"02";
            when "00" & x"852" => data <= x"a2";
            when "00" & x"853" => data <= x"02";
            when "00" & x"854" => data <= x"20";
            when "00" & x"855" => data <= x"60";
            when "00" & x"856" => data <= x"88";
            when "00" & x"857" => data <= x"9d";
            when "00" & x"858" => data <= x"cb";
            when "00" & x"859" => data <= x"10";
            when "00" & x"85a" => data <= x"a5";
            when "00" & x"85b" => data <= x"ce";
            when "00" & x"85c" => data <= x"9d";
            when "00" & x"85d" => data <= x"ca";
            when "00" & x"85e" => data <= x"10";
            when "00" & x"85f" => data <= x"60";
            when "00" & x"860" => data <= x"a9";
            when "00" & x"861" => data <= x"24";
            when "00" & x"862" => data <= x"85";
            when "00" & x"863" => data <= x"ce";
            when "00" & x"864" => data <= x"20";
            when "00" & x"865" => data <= x"bf";
            when "00" & x"866" => data <= x"86";
            when "00" & x"867" => data <= x"d0";
            when "00" & x"868" => data <= x"07";
            when "00" & x"869" => data <= x"a9";
            when "00" & x"86a" => data <= x"00";
            when "00" & x"86b" => data <= x"20";
            when "00" & x"86c" => data <= x"7e";
            when "00" & x"86d" => data <= x"87";
            when "00" & x"86e" => data <= x"f0";
            when "00" & x"86f" => data <= x"30";
            when "00" & x"870" => data <= x"ad";
            when "00" & x"871" => data <= x"cb";
            when "00" & x"872" => data <= x"10";
            when "00" & x"873" => data <= x"20";
            when "00" & x"874" => data <= x"7e";
            when "00" & x"875" => data <= x"87";
            when "00" & x"876" => data <= x"20";
            when "00" & x"877" => data <= x"c5";
            when "00" & x"878" => data <= x"ff";
            when "00" & x"879" => data <= x"b0";
            when "00" & x"87a" => data <= x"10";
            when "00" & x"87b" => data <= x"c9";
            when "00" & x"87c" => data <= x"3a";
            when "00" & x"87d" => data <= x"d0";
            when "00" & x"87e" => data <= x"1a";
            when "00" & x"87f" => data <= x"20";
            when "00" & x"880" => data <= x"5d";
            when "00" & x"881" => data <= x"83";
            when "00" & x"882" => data <= x"20";
            when "00" & x"883" => data <= x"c5";
            when "00" & x"884" => data <= x"ff";
            when "00" & x"885" => data <= x"b0";
            when "00" & x"886" => data <= x"19";
            when "00" & x"887" => data <= x"c9";
            when "00" & x"888" => data <= x"2e";
            when "00" & x"889" => data <= x"f0";
            when "00" & x"88a" => data <= x"eb";
            when "00" & x"88b" => data <= x"20";
            when "00" & x"88c" => data <= x"22";
            when "00" & x"88d" => data <= x"80";
            when "00" & x"88e" => data <= x"ce";
            when "00" & x"88f" => data <= x"64";
            when "00" & x"890" => data <= x"69";
            when "00" & x"891" => data <= x"72";
            when "00" & x"892" => data <= x"65";
            when "00" & x"893" => data <= x"63";
            when "00" & x"894" => data <= x"74";
            when "00" & x"895" => data <= x"6f";
            when "00" & x"896" => data <= x"72";
            when "00" & x"897" => data <= x"79";
            when "00" & x"898" => data <= x"00";
            when "00" & x"899" => data <= x"85";
            when "00" & x"89a" => data <= x"ce";
            when "00" & x"89b" => data <= x"20";
            when "00" & x"89c" => data <= x"c5";
            when "00" & x"89d" => data <= x"ff";
            when "00" & x"89e" => data <= x"90";
            when "00" & x"89f" => data <= x"eb";
            when "00" & x"8a0" => data <= x"a5";
            when "00" & x"8a1" => data <= x"cf";
            when "00" & x"8a2" => data <= x"60";
            when "00" & x"8a3" => data <= x"20";
            when "00" & x"8a4" => data <= x"01";
            when "00" & x"8a5" => data <= x"9a";
            when "00" & x"8a6" => data <= x"20";
            when "00" & x"8a7" => data <= x"4d";
            when "00" & x"8a8" => data <= x"83";
            when "00" & x"8a9" => data <= x"20";
            when "00" & x"8aa" => data <= x"47";
            when "00" & x"8ab" => data <= x"83";
            when "00" & x"8ac" => data <= x"4c";
            when "00" & x"8ad" => data <= x"ce";
            when "00" & x"8ae" => data <= x"b2";
            when "00" & x"8af" => data <= x"00";
            when "00" & x"8b0" => data <= x"20";
            when "00" & x"8b1" => data <= x"c6";
            when "00" & x"8b2" => data <= x"88";
            when "00" & x"8b3" => data <= x"ca";
            when "00" & x"8b4" => data <= x"10";
            when "00" & x"8b5" => data <= x"fa";
            when "00" & x"8b6" => data <= x"e8";
            when "00" & x"8b7" => data <= x"20";
            when "00" & x"8b8" => data <= x"c5";
            when "00" & x"8b9" => data <= x"ff";
            when "00" & x"8ba" => data <= x"b0";
            when "00" & x"8bb" => data <= x"07";
            when "00" & x"8bc" => data <= x"20";
            when "00" & x"8bd" => data <= x"c6";
            when "00" & x"8be" => data <= x"88";
            when "00" & x"8bf" => data <= x"e0";
            when "00" & x"8c0" => data <= x"0b";
            when "00" & x"8c1" => data <= x"90";
            when "00" & x"8c2" => data <= x"f3";
            when "00" & x"8c3" => data <= x"4c";
            when "00" & x"8c4" => data <= x"b4";
            when "00" & x"8c5" => data <= x"8a";
            when "00" & x"8c6" => data <= x"e0";
            when "00" & x"8c7" => data <= x"08";
            when "00" & x"8c8" => data <= x"90";
            when "00" & x"8c9" => data <= x"04";
            when "00" & x"8ca" => data <= x"9d";
            when "00" & x"8cb" => data <= x"f8";
            when "00" & x"8cc" => data <= x"0e";
            when "00" & x"8cd" => data <= x"60";
            when "00" & x"8ce" => data <= x"9d";
            when "00" & x"8cf" => data <= x"00";
            when "00" & x"8d0" => data <= x"0e";
            when "00" & x"8d1" => data <= x"60";
            when "00" & x"8d2" => data <= x"20";
            when "00" & x"8d3" => data <= x"5e";
            when "00" & x"8d4" => data <= x"82";
            when "00" & x"8d5" => data <= x"20";
            when "00" & x"8d6" => data <= x"01";
            when "00" & x"8d7" => data <= x"9a";
            when "00" & x"8d8" => data <= x"20";
            when "00" & x"8d9" => data <= x"fe";
            when "00" & x"8da" => data <= x"80";
            when "00" & x"8db" => data <= x"a2";
            when "00" & x"8dc" => data <= x"00";
            when "00" & x"8dd" => data <= x"20";
            when "00" & x"8de" => data <= x"bf";
            when "00" & x"8df" => data <= x"86";
            when "00" & x"8e0" => data <= x"d0";
            when "00" & x"8e1" => data <= x"23";
            when "00" & x"8e2" => data <= x"86";
            when "00" & x"8e3" => data <= x"aa";
            when "00" & x"8e4" => data <= x"20";
            when "00" & x"8e5" => data <= x"96";
            when "00" & x"8e6" => data <= x"82";
            when "00" & x"8e7" => data <= x"b0";
            when "00" & x"8e8" => data <= x"03";
            when "00" & x"8e9" => data <= x"4c";
            when "00" & x"8ea" => data <= x"76";
            when "00" & x"8eb" => data <= x"82";
            when "00" & x"8ec" => data <= x"20";
            when "00" & x"8ed" => data <= x"4f";
            when "00" & x"8ee" => data <= x"98";
            when "00" & x"8ef" => data <= x"b9";
            when "00" & x"8f0" => data <= x"0f";
            when "00" & x"8f1" => data <= x"0e";
            when "00" & x"8f2" => data <= x"29";
            when "00" & x"8f3" => data <= x"7f";
            when "00" & x"8f4" => data <= x"05";
            when "00" & x"8f5" => data <= x"aa";
            when "00" & x"8f6" => data <= x"99";
            when "00" & x"8f7" => data <= x"0f";
            when "00" & x"8f8" => data <= x"0e";
            when "00" & x"8f9" => data <= x"20";
            when "00" & x"8fa" => data <= x"fc";
            when "00" & x"8fb" => data <= x"82";
            when "00" & x"8fc" => data <= x"20";
            when "00" & x"8fd" => data <= x"9d";
            when "00" & x"8fe" => data <= x"82";
            when "00" & x"8ff" => data <= x"b0";
            when "00" & x"900" => data <= x"eb";
            when "00" & x"901" => data <= x"90";
            when "00" & x"902" => data <= x"c0";
            when "00" & x"903" => data <= x"a2";
            when "00" & x"904" => data <= x"80";
            when "00" & x"905" => data <= x"20";
            when "00" & x"906" => data <= x"c5";
            when "00" & x"907" => data <= x"ff";
            when "00" & x"908" => data <= x"b0";
            when "00" & x"909" => data <= x"d8";
            when "00" & x"90a" => data <= x"c9";
            when "00" & x"90b" => data <= x"4c";
            when "00" & x"90c" => data <= x"f0";
            when "00" & x"90d" => data <= x"f5";
            when "00" & x"90e" => data <= x"20";
            when "00" & x"90f" => data <= x"22";
            when "00" & x"910" => data <= x"80";
            when "00" & x"911" => data <= x"cf";
            when "00" & x"912" => data <= x"61";
            when "00" & x"913" => data <= x"74";
            when "00" & x"914" => data <= x"74";
            when "00" & x"915" => data <= x"72";
            when "00" & x"916" => data <= x"69";
            when "00" & x"917" => data <= x"62";
            when "00" & x"918" => data <= x"75";
            when "00" & x"919" => data <= x"74";
            when "00" & x"91a" => data <= x"65";
            when "00" & x"91b" => data <= x"00";
            when "00" & x"91c" => data <= x"20";
            when "00" & x"91d" => data <= x"e1";
            when "00" & x"91e" => data <= x"83";
            when "00" & x"91f" => data <= x"8a";
            when "00" & x"920" => data <= x"c9";
            when "00" & x"921" => data <= x"04";
            when "00" & x"922" => data <= x"f0";
            when "00" & x"923" => data <= x"1a";
            when "00" & x"924" => data <= x"c9";
            when "00" & x"925" => data <= x"02";
            when "00" & x"926" => data <= x"90";
            when "00" & x"927" => data <= x"0b";
            when "00" & x"928" => data <= x"20";
            when "00" & x"929" => data <= x"22";
            when "00" & x"92a" => data <= x"80";
            when "00" & x"92b" => data <= x"cb";
            when "00" & x"92c" => data <= x"6f";
            when "00" & x"92d" => data <= x"70";
            when "00" & x"92e" => data <= x"74";
            when "00" & x"92f" => data <= x"69";
            when "00" & x"930" => data <= x"6f";
            when "00" & x"931" => data <= x"6e";
            when "00" & x"932" => data <= x"00";
            when "00" & x"933" => data <= x"a2";
            when "00" & x"934" => data <= x"ff";
            when "00" & x"935" => data <= x"98";
            when "00" & x"936" => data <= x"f0";
            when "00" & x"937" => data <= x"02";
            when "00" & x"938" => data <= x"a2";
            when "00" & x"939" => data <= x"00";
            when "00" & x"93a" => data <= x"8e";
            when "00" & x"93b" => data <= x"c7";
            when "00" & x"93c" => data <= x"10";
            when "00" & x"93d" => data <= x"60";
            when "00" & x"93e" => data <= x"98";
            when "00" & x"93f" => data <= x"48";
            when "00" & x"940" => data <= x"20";
            when "00" & x"941" => data <= x"4d";
            when "00" & x"942" => data <= x"83";
            when "00" & x"943" => data <= x"20";
            when "00" & x"944" => data <= x"41";
            when "00" & x"945" => data <= x"af";
            when "00" & x"946" => data <= x"68";
            when "00" & x"947" => data <= x"20";
            when "00" & x"948" => data <= x"0b";
            when "00" & x"949" => data <= x"82";
            when "00" & x"94a" => data <= x"4d";
            when "00" & x"94b" => data <= x"06";
            when "00" & x"94c" => data <= x"0f";
            when "00" & x"94d" => data <= x"29";
            when "00" & x"94e" => data <= x"30";
            when "00" & x"94f" => data <= x"4d";
            when "00" & x"950" => data <= x"06";
            when "00" & x"951" => data <= x"0f";
            when "00" & x"952" => data <= x"8d";
            when "00" & x"953" => data <= x"06";
            when "00" & x"954" => data <= x"0f";
            when "00" & x"955" => data <= x"4c";
            when "00" & x"956" => data <= x"b4";
            when "00" & x"957" => data <= x"8a";
            when "00" & x"958" => data <= x"20";
            when "00" & x"959" => data <= x"18";
            when "00" & x"95a" => data <= x"80";
            when "00" & x"95b" => data <= x"c6";
            when "00" & x"95c" => data <= x"66";
            when "00" & x"95d" => data <= x"75";
            when "00" & x"95e" => data <= x"6c";
            when "00" & x"95f" => data <= x"6c";
            when "00" & x"960" => data <= x"00";
            when "00" & x"961" => data <= x"20";
            when "00" & x"962" => data <= x"06";
            when "00" & x"963" => data <= x"81";
            when "00" & x"964" => data <= x"20";
            when "00" & x"965" => data <= x"96";
            when "00" & x"966" => data <= x"82";
            when "00" & x"967" => data <= x"90";
            when "00" & x"968" => data <= x"03";
            when "00" & x"969" => data <= x"20";
            when "00" & x"96a" => data <= x"d1";
            when "00" & x"96b" => data <= x"82";
            when "00" & x"96c" => data <= x"a5";
            when "00" & x"96d" => data <= x"c2";
            when "00" & x"96e" => data <= x"48";
            when "00" & x"96f" => data <= x"a5";
            when "00" & x"970" => data <= x"c3";
            when "00" & x"971" => data <= x"48";
            when "00" & x"972" => data <= x"38";
            when "00" & x"973" => data <= x"a5";
            when "00" & x"974" => data <= x"c4";
            when "00" & x"975" => data <= x"e5";
            when "00" & x"976" => data <= x"c2";
            when "00" & x"977" => data <= x"85";
            when "00" & x"978" => data <= x"c2";
            when "00" & x"979" => data <= x"a5";
            when "00" & x"97a" => data <= x"c5";
            when "00" & x"97b" => data <= x"e5";
            when "00" & x"97c" => data <= x"c3";
            when "00" & x"97d" => data <= x"85";
            when "00" & x"97e" => data <= x"c3";
            when "00" & x"97f" => data <= x"ad";
            when "00" & x"980" => data <= x"7a";
            when "00" & x"981" => data <= x"10";
            when "00" & x"982" => data <= x"ed";
            when "00" & x"983" => data <= x"78";
            when "00" & x"984" => data <= x"10";
            when "00" & x"985" => data <= x"85";
            when "00" & x"986" => data <= x"c6";
            when "00" & x"987" => data <= x"20";
            when "00" & x"988" => data <= x"9d";
            when "00" & x"989" => data <= x"89";
            when "00" & x"98a" => data <= x"ad";
            when "00" & x"98b" => data <= x"79";
            when "00" & x"98c" => data <= x"10";
            when "00" & x"98d" => data <= x"8d";
            when "00" & x"98e" => data <= x"75";
            when "00" & x"98f" => data <= x"10";
            when "00" & x"990" => data <= x"ad";
            when "00" & x"991" => data <= x"78";
            when "00" & x"992" => data <= x"10";
            when "00" & x"993" => data <= x"8d";
            when "00" & x"994" => data <= x"74";
            when "00" & x"995" => data <= x"10";
            when "00" & x"996" => data <= x"68";
            when "00" & x"997" => data <= x"85";
            when "00" & x"998" => data <= x"bf";
            when "00" & x"999" => data <= x"68";
            when "00" & x"99a" => data <= x"85";
            when "00" & x"99b" => data <= x"be";
            when "00" & x"99c" => data <= x"60";
            when "00" & x"99d" => data <= x"a9";
            when "00" & x"99e" => data <= x"00";
            when "00" & x"99f" => data <= x"85";
            when "00" & x"9a0" => data <= x"c4";
            when "00" & x"9a1" => data <= x"a9";
            when "00" & x"9a2" => data <= x"02";
            when "00" & x"9a3" => data <= x"85";
            when "00" & x"9a4" => data <= x"c5";
            when "00" & x"9a5" => data <= x"ac";
            when "00" & x"9a6" => data <= x"05";
            when "00" & x"9a7" => data <= x"0f";
            when "00" & x"9a8" => data <= x"f0";
            when "00" & x"9a9" => data <= x"2d";
            when "00" & x"9aa" => data <= x"c0";
            when "00" & x"9ab" => data <= x"f8";
            when "00" & x"9ac" => data <= x"b0";
            when "00" & x"9ad" => data <= x"56";
            when "00" & x"9ae" => data <= x"20";
            when "00" & x"9af" => data <= x"9e";
            when "00" & x"9b0" => data <= x"85";
            when "00" & x"9b1" => data <= x"4c";
            when "00" & x"9b2" => data <= x"bc";
            when "00" & x"9b3" => data <= x"89";
            when "00" & x"9b4" => data <= x"f0";
            when "00" & x"9b5" => data <= x"a2";
            when "00" & x"9b6" => data <= x"20";
            when "00" & x"9b7" => data <= x"19";
            when "00" & x"9b8" => data <= x"82";
            when "00" & x"9b9" => data <= x"20";
            when "00" & x"9ba" => data <= x"7f";
            when "00" & x"9bb" => data <= x"85";
            when "00" & x"9bc" => data <= x"98";
            when "00" & x"9bd" => data <= x"90";
            when "00" & x"9be" => data <= x"f5";
            when "00" & x"9bf" => data <= x"84";
            when "00" & x"9c0" => data <= x"b0";
            when "00" & x"9c1" => data <= x"ac";
            when "00" & x"9c2" => data <= x"05";
            when "00" & x"9c3" => data <= x"0f";
            when "00" & x"9c4" => data <= x"c4";
            when "00" & x"9c5" => data <= x"b0";
            when "00" & x"9c6" => data <= x"f0";
            when "00" & x"9c7" => data <= x"0f";
            when "00" & x"9c8" => data <= x"b9";
            when "00" & x"9c9" => data <= x"07";
            when "00" & x"9ca" => data <= x"0e";
            when "00" & x"9cb" => data <= x"99";
            when "00" & x"9cc" => data <= x"0f";
            when "00" & x"9cd" => data <= x"0e";
            when "00" & x"9ce" => data <= x"b9";
            when "00" & x"9cf" => data <= x"07";
            when "00" & x"9d0" => data <= x"0f";
            when "00" & x"9d1" => data <= x"99";
            when "00" & x"9d2" => data <= x"0f";
            when "00" & x"9d3" => data <= x"0f";
            when "00" & x"9d4" => data <= x"88";
            when "00" & x"9d5" => data <= x"b0";
            when "00" & x"9d6" => data <= x"ed";
            when "00" & x"9d7" => data <= x"a2";
            when "00" & x"9d8" => data <= x"00";
            when "00" & x"9d9" => data <= x"20";
            when "00" & x"9da" => data <= x"17";
            when "00" & x"9db" => data <= x"8a";
            when "00" & x"9dc" => data <= x"b5";
            when "00" & x"9dd" => data <= x"c7";
            when "00" & x"9de" => data <= x"99";
            when "00" & x"9df" => data <= x"08";
            when "00" & x"9e0" => data <= x"0e";
            when "00" & x"9e1" => data <= x"c8";
            when "00" & x"9e2" => data <= x"e8";
            when "00" & x"9e3" => data <= x"e0";
            when "00" & x"9e4" => data <= x"08";
            when "00" & x"9e5" => data <= x"d0";
            when "00" & x"9e6" => data <= x"f5";
            when "00" & x"9e7" => data <= x"b5";
            when "00" & x"9e8" => data <= x"bd";
            when "00" & x"9e9" => data <= x"88";
            when "00" & x"9ea" => data <= x"99";
            when "00" & x"9eb" => data <= x"08";
            when "00" & x"9ec" => data <= x"0f";
            when "00" & x"9ed" => data <= x"ca";
            when "00" & x"9ee" => data <= x"d0";
            when "00" & x"9ef" => data <= x"f7";
            when "00" & x"9f0" => data <= x"20";
            when "00" & x"9f1" => data <= x"fc";
            when "00" & x"9f2" => data <= x"82";
            when "00" & x"9f3" => data <= x"98";
            when "00" & x"9f4" => data <= x"48";
            when "00" & x"9f5" => data <= x"ac";
            when "00" & x"9f6" => data <= x"05";
            when "00" & x"9f7" => data <= x"0f";
            when "00" & x"9f8" => data <= x"20";
            when "00" & x"9f9" => data <= x"10";
            when "00" & x"9fa" => data <= x"82";
            when "00" & x"9fb" => data <= x"8c";
            when "00" & x"9fc" => data <= x"05";
            when "00" & x"9fd" => data <= x"0f";
            when "00" & x"9fe" => data <= x"20";
            when "00" & x"9ff" => data <= x"b4";
            when "00" & x"a00" => data <= x"8a";
            when "00" & x"a01" => data <= x"68";
            when "00" & x"a02" => data <= x"a8";
            when "00" & x"a03" => data <= x"60";
            when "00" & x"a04" => data <= x"20";
            when "00" & x"a05" => data <= x"33";
            when "00" & x"a06" => data <= x"80";
            when "00" & x"a07" => data <= x"be";
            when "00" & x"a08" => data <= x"43";
            when "00" & x"a09" => data <= x"61";
            when "00" & x"a0a" => data <= x"74";
            when "00" & x"a0b" => data <= x"61";
            when "00" & x"a0c" => data <= x"6c";
            when "00" & x"a0d" => data <= x"6f";
            when "00" & x"a0e" => data <= x"67";
            when "00" & x"a0f" => data <= x"75";
            when "00" & x"a10" => data <= x"65";
            when "00" & x"a11" => data <= x"20";
            when "00" & x"a12" => data <= x"66";
            when "00" & x"a13" => data <= x"75";
            when "00" & x"a14" => data <= x"6c";
            when "00" & x"a15" => data <= x"6c";
            when "00" & x"a16" => data <= x"00";
            when "00" & x"a17" => data <= x"ad";
            when "00" & x"a18" => data <= x"76";
            when "00" & x"a19" => data <= x"10";
            when "00" & x"a1a" => data <= x"29";
            when "00" & x"a1b" => data <= x"03";
            when "00" & x"a1c" => data <= x"0a";
            when "00" & x"a1d" => data <= x"0a";
            when "00" & x"a1e" => data <= x"45";
            when "00" & x"a1f" => data <= x"c6";
            when "00" & x"a20" => data <= x"29";
            when "00" & x"a21" => data <= x"fc";
            when "00" & x"a22" => data <= x"45";
            when "00" & x"a23" => data <= x"c6";
            when "00" & x"a24" => data <= x"0a";
            when "00" & x"a25" => data <= x"0a";
            when "00" & x"a26" => data <= x"4d";
            when "00" & x"a27" => data <= x"74";
            when "00" & x"a28" => data <= x"10";
            when "00" & x"a29" => data <= x"29";
            when "00" & x"a2a" => data <= x"fc";
            when "00" & x"a2b" => data <= x"4d";
            when "00" & x"a2c" => data <= x"74";
            when "00" & x"a2d" => data <= x"10";
            when "00" & x"a2e" => data <= x"0a";
            when "00" & x"a2f" => data <= x"0a";
            when "00" & x"a30" => data <= x"45";
            when "00" & x"a31" => data <= x"c4";
            when "00" & x"a32" => data <= x"29";
            when "00" & x"a33" => data <= x"fc";
            when "00" & x"a34" => data <= x"45";
            when "00" & x"a35" => data <= x"c4";
            when "00" & x"a36" => data <= x"85";
            when "00" & x"a37" => data <= x"c4";
            when "00" & x"a38" => data <= x"60";
            when "00" & x"a39" => data <= x"a9";
            when "00" & x"a3a" => data <= x"01";
            when "00" & x"a3b" => data <= x"8d";
            when "00" & x"a3c" => data <= x"c8";
            when "00" & x"a3d" => data <= x"10";
            when "00" & x"a3e" => data <= x"60";
            when "00" & x"a3f" => data <= x"a9";
            when "00" & x"a40" => data <= x"00";
            when "00" & x"a41" => data <= x"8d";
            when "00" & x"a42" => data <= x"75";
            when "00" & x"a43" => data <= x"10";
            when "00" & x"a44" => data <= x"a5";
            when "00" & x"a45" => data <= x"c4";
            when "00" & x"a46" => data <= x"20";
            when "00" & x"a47" => data <= x"ff";
            when "00" & x"a48" => data <= x"81";
            when "00" & x"a49" => data <= x"c9";
            when "00" & x"a4a" => data <= x"03";
            when "00" & x"a4b" => data <= x"d0";
            when "00" & x"a4c" => data <= x"05";
            when "00" & x"a4d" => data <= x"a9";
            when "00" & x"a4e" => data <= x"ff";
            when "00" & x"a4f" => data <= x"8d";
            when "00" & x"a50" => data <= x"75";
            when "00" & x"a51" => data <= x"10";
            when "00" & x"a52" => data <= x"8d";
            when "00" & x"a53" => data <= x"74";
            when "00" & x"a54" => data <= x"10";
            when "00" & x"a55" => data <= x"60";
            when "00" & x"a56" => data <= x"a9";
            when "00" & x"a57" => data <= x"00";
            when "00" & x"a58" => data <= x"8d";
            when "00" & x"a59" => data <= x"77";
            when "00" & x"a5a" => data <= x"10";
            when "00" & x"a5b" => data <= x"a5";
            when "00" & x"a5c" => data <= x"c4";
            when "00" & x"a5d" => data <= x"20";
            when "00" & x"a5e" => data <= x"fb";
            when "00" & x"a5f" => data <= x"81";
            when "00" & x"a60" => data <= x"c9";
            when "00" & x"a61" => data <= x"03";
            when "00" & x"a62" => data <= x"d0";
            when "00" & x"a63" => data <= x"05";
            when "00" & x"a64" => data <= x"a9";
            when "00" & x"a65" => data <= x"ff";
            when "00" & x"a66" => data <= x"8d";
            when "00" & x"a67" => data <= x"77";
            when "00" & x"a68" => data <= x"10";
            when "00" & x"a69" => data <= x"8d";
            when "00" & x"a6a" => data <= x"76";
            when "00" & x"a6b" => data <= x"10";
            when "00" & x"a6c" => data <= x"60";
            when "00" & x"a6d" => data <= x"20";
            when "00" & x"a6e" => data <= x"62";
            when "00" & x"a6f" => data <= x"82";
            when "00" & x"a70" => data <= x"20";
            when "00" & x"a71" => data <= x"bf";
            when "00" & x"a72" => data <= x"86";
            when "00" & x"a73" => data <= x"d0";
            when "00" & x"a74" => data <= x"03";
            when "00" & x"a75" => data <= x"4c";
            when "00" & x"a76" => data <= x"06";
            when "00" & x"a77" => data <= x"9a";
            when "00" & x"a78" => data <= x"20";
            when "00" & x"a79" => data <= x"fe";
            when "00" & x"a7a" => data <= x"80";
            when "00" & x"a7b" => data <= x"98";
            when "00" & x"a7c" => data <= x"48";
            when "00" & x"a7d" => data <= x"20";
            when "00" & x"a7e" => data <= x"96";
            when "00" & x"a7f" => data <= x"82";
            when "00" & x"a80" => data <= x"b0";
            when "00" & x"a81" => data <= x"03";
            when "00" & x"a82" => data <= x"4c";
            when "00" & x"a83" => data <= x"76";
            when "00" & x"a84" => data <= x"82";
            when "00" & x"a85" => data <= x"20";
            when "00" & x"a86" => data <= x"4c";
            when "00" & x"a87" => data <= x"98";
            when "00" & x"a88" => data <= x"84";
            when "00" & x"a89" => data <= x"b3";
            when "00" & x"a8a" => data <= x"68";
            when "00" & x"a8b" => data <= x"a8";
            when "00" & x"a8c" => data <= x"20";
            when "00" & x"a8d" => data <= x"bf";
            when "00" & x"a8e" => data <= x"86";
            when "00" & x"a8f" => data <= x"f0";
            when "00" & x"a90" => data <= x"e4";
            when "00" & x"a91" => data <= x"20";
            when "00" & x"a92" => data <= x"fe";
            when "00" & x"a93" => data <= x"80";
            when "00" & x"a94" => data <= x"20";
            when "00" & x"a95" => data <= x"96";
            when "00" & x"a96" => data <= x"82";
            when "00" & x"a97" => data <= x"90";
            when "00" & x"a98" => data <= x"0b";
            when "00" & x"a99" => data <= x"20";
            when "00" & x"a9a" => data <= x"2b";
            when "00" & x"a9b" => data <= x"80";
            when "00" & x"a9c" => data <= x"c4";
            when "00" & x"a9d" => data <= x"65";
            when "00" & x"a9e" => data <= x"78";
            when "00" & x"a9f" => data <= x"69";
            when "00" & x"aa0" => data <= x"73";
            when "00" & x"aa1" => data <= x"74";
            when "00" & x"aa2" => data <= x"73";
            when "00" & x"aa3" => data <= x"00";
            when "00" & x"aa4" => data <= x"a4";
            when "00" & x"aa5" => data <= x"b3";
            when "00" & x"aa6" => data <= x"20";
            when "00" & x"aa7" => data <= x"10";
            when "00" & x"aa8" => data <= x"82";
            when "00" & x"aa9" => data <= x"a2";
            when "00" & x"aaa" => data <= x"07";
            when "00" & x"aab" => data <= x"b5";
            when "00" & x"aac" => data <= x"c7";
            when "00" & x"aad" => data <= x"99";
            when "00" & x"aae" => data <= x"07";
            when "00" & x"aaf" => data <= x"0e";
            when "00" & x"ab0" => data <= x"88";
            when "00" & x"ab1" => data <= x"ca";
            when "00" & x"ab2" => data <= x"10";
            when "00" & x"ab3" => data <= x"f7";
            when "00" & x"ab4" => data <= x"18";
            when "00" & x"ab5" => data <= x"f8";
            when "00" & x"ab6" => data <= x"ad";
            when "00" & x"ab7" => data <= x"04";
            when "00" & x"ab8" => data <= x"0f";
            when "00" & x"ab9" => data <= x"69";
            when "00" & x"aba" => data <= x"01";
            when "00" & x"abb" => data <= x"d8";
            when "00" & x"abc" => data <= x"8d";
            when "00" & x"abd" => data <= x"04";
            when "00" & x"abe" => data <= x"0f";
            when "00" & x"abf" => data <= x"4c";
            when "00" & x"ac0" => data <= x"55";
            when "00" & x"ac1" => data <= x"af";
            when "00" & x"ac2" => data <= x"a9";
            when "00" & x"ac3" => data <= x"ff";
            when "00" & x"ac4" => data <= x"20";
            when "00" & x"ac5" => data <= x"9e";
            when "00" & x"ac6" => data <= x"06";
            when "00" & x"ac7" => data <= x"ad";
            when "00" & x"ac8" => data <= x"e3";
            when "00" & x"ac9" => data <= x"fe";
            when "00" & x"aca" => data <= x"a9";
            when "00" & x"acb" => data <= x"00";
            when "00" & x"acc" => data <= x"20";
            when "00" & x"acd" => data <= x"95";
            when "00" & x"ace" => data <= x"06";
            when "00" & x"acf" => data <= x"a8";
            when "00" & x"ad0" => data <= x"b1";
            when "00" & x"ad1" => data <= x"fd";
            when "00" & x"ad2" => data <= x"20";
            when "00" & x"ad3" => data <= x"95";
            when "00" & x"ad4" => data <= x"06";
            when "00" & x"ad5" => data <= x"c8";
            when "00" & x"ad6" => data <= x"b1";
            when "00" & x"ad7" => data <= x"fd";
            when "00" & x"ad8" => data <= x"20";
            when "00" & x"ad9" => data <= x"95";
            when "00" & x"ada" => data <= x"06";
            when "00" & x"adb" => data <= x"aa";
            when "00" & x"adc" => data <= x"d0";
            when "00" & x"add" => data <= x"f7";
            when "00" & x"ade" => data <= x"a2";
            when "00" & x"adf" => data <= x"ff";
            when "00" & x"ae0" => data <= x"9a";
            when "00" & x"ae1" => data <= x"58";
            when "00" & x"ae2" => data <= x"2c";
            when "00" & x"ae3" => data <= x"e0";
            when "00" & x"ae4" => data <= x"fe";
            when "00" & x"ae5" => data <= x"10";
            when "00" & x"ae6" => data <= x"06";
            when "00" & x"ae7" => data <= x"ad";
            when "00" & x"ae8" => data <= x"e1";
            when "00" & x"ae9" => data <= x"fe";
            when "00" & x"aea" => data <= x"20";
            when "00" & x"aeb" => data <= x"ee";
            when "00" & x"aec" => data <= x"ff";
            when "00" & x"aed" => data <= x"2c";
            when "00" & x"aee" => data <= x"e2";
            when "00" & x"aef" => data <= x"fe";
            when "00" & x"af0" => data <= x"10";
            when "00" & x"af1" => data <= x"f0";
            when "00" & x"af2" => data <= x"2c";
            when "00" & x"af3" => data <= x"e0";
            when "00" & x"af4" => data <= x"fe";
            when "00" & x"af5" => data <= x"30";
            when "00" & x"af6" => data <= x"f0";
            when "00" & x"af7" => data <= x"ae";
            when "00" & x"af8" => data <= x"e3";
            when "00" & x"af9" => data <= x"fe";
            when "00" & x"afa" => data <= x"86";
            when "00" & x"afb" => data <= x"51";
            when "00" & x"afc" => data <= x"6c";
            when "00" & x"afd" => data <= x"00";
            when "00" & x"afe" => data <= x"05";
            when "00" & x"aff" => data <= x"00";
            when "00" & x"b00" => data <= x"80";
            when "00" & x"b01" => data <= x"00";
            when "00" & x"b02" => data <= x"00";
            when "00" & x"b03" => data <= x"4c";
            when "00" & x"b04" => data <= x"84";
            when "00" & x"b05" => data <= x"04";
            when "00" & x"b06" => data <= x"4c";
            when "00" & x"b07" => data <= x"a7";
            when "00" & x"b08" => data <= x"06";
            when "00" & x"b09" => data <= x"c9";
            when "00" & x"b0a" => data <= x"80";
            when "00" & x"b0b" => data <= x"90";
            when "00" & x"b0c" => data <= x"2b";
            when "00" & x"b0d" => data <= x"c9";
            when "00" & x"b0e" => data <= x"c0";
            when "00" & x"b0f" => data <= x"b0";
            when "00" & x"b10" => data <= x"1a";
            when "00" & x"b11" => data <= x"09";
            when "00" & x"b12" => data <= x"40";
            when "00" & x"b13" => data <= x"c5";
            when "00" & x"b14" => data <= x"15";
            when "00" & x"b15" => data <= x"d0";
            when "00" & x"b16" => data <= x"20";
            when "00" & x"b17" => data <= x"08";
            when "00" & x"b18" => data <= x"78";
            when "00" & x"b19" => data <= x"a9";
            when "00" & x"b1a" => data <= x"05";
            when "00" & x"b1b" => data <= x"20";
            when "00" & x"b1c" => data <= x"9e";
            when "00" & x"b1d" => data <= x"06";
            when "00" & x"b1e" => data <= x"a5";
            when "00" & x"b1f" => data <= x"15";
            when "00" & x"b20" => data <= x"20";
            when "00" & x"b21" => data <= x"9e";
            when "00" & x"b22" => data <= x"06";
            when "00" & x"b23" => data <= x"28";
            when "00" & x"b24" => data <= x"a9";
            when "00" & x"b25" => data <= x"80";
            when "00" & x"b26" => data <= x"85";
            when "00" & x"b27" => data <= x"15";
            when "00" & x"b28" => data <= x"85";
            when "00" & x"b29" => data <= x"14";
            when "00" & x"b2a" => data <= x"60";
            when "00" & x"b2b" => data <= x"06";
            when "00" & x"b2c" => data <= x"14";
            when "00" & x"b2d" => data <= x"b0";
            when "00" & x"b2e" => data <= x"06";
            when "00" & x"b2f" => data <= x"c5";
            when "00" & x"b30" => data <= x"15";
            when "00" & x"b31" => data <= x"f0";
            when "00" & x"b32" => data <= x"04";
            when "00" & x"b33" => data <= x"18";
            when "00" & x"b34" => data <= x"60";
            when "00" & x"b35" => data <= x"85";
            when "00" & x"b36" => data <= x"15";
            when "00" & x"b37" => data <= x"60";
            when "00" & x"b38" => data <= x"08";
            when "00" & x"b39" => data <= x"78";
            when "00" & x"b3a" => data <= x"84";
            when "00" & x"b3b" => data <= x"13";
            when "00" & x"b3c" => data <= x"86";
            when "00" & x"b3d" => data <= x"12";
            when "00" & x"b3e" => data <= x"20";
            when "00" & x"b3f" => data <= x"9e";
            when "00" & x"b40" => data <= x"06";
            when "00" & x"b41" => data <= x"aa";
            when "00" & x"b42" => data <= x"a0";
            when "00" & x"b43" => data <= x"03";
            when "00" & x"b44" => data <= x"a5";
            when "00" & x"b45" => data <= x"15";
            when "00" & x"b46" => data <= x"20";
            when "00" & x"b47" => data <= x"9e";
            when "00" & x"b48" => data <= x"06";
            when "00" & x"b49" => data <= x"b1";
            when "00" & x"b4a" => data <= x"12";
            when "00" & x"b4b" => data <= x"20";
            when "00" & x"b4c" => data <= x"9e";
            when "00" & x"b4d" => data <= x"06";
            when "00" & x"b4e" => data <= x"88";
            when "00" & x"b4f" => data <= x"10";
            when "00" & x"b50" => data <= x"f8";
            when "00" & x"b51" => data <= x"a0";
            when "00" & x"b52" => data <= x"18";
            when "00" & x"b53" => data <= x"8c";
            when "00" & x"b54" => data <= x"e0";
            when "00" & x"b55" => data <= x"fe";
            when "00" & x"b56" => data <= x"bd";
            when "00" & x"b57" => data <= x"18";
            when "00" & x"b58" => data <= x"05";
            when "00" & x"b59" => data <= x"8d";
            when "00" & x"b5a" => data <= x"e0";
            when "00" & x"b5b" => data <= x"fe";
            when "00" & x"b5c" => data <= x"4a";
            when "00" & x"b5d" => data <= x"4a";
            when "00" & x"b5e" => data <= x"90";
            when "00" & x"b5f" => data <= x"06";
            when "00" & x"b60" => data <= x"2c";
            when "00" & x"b61" => data <= x"e5";
            when "00" & x"b62" => data <= x"fe";
            when "00" & x"b63" => data <= x"2c";
            when "00" & x"b64" => data <= x"e5";
            when "00" & x"b65" => data <= x"fe";
            when "00" & x"b66" => data <= x"20";
            when "00" & x"b67" => data <= x"9e";
            when "00" & x"b68" => data <= x"06";
            when "00" & x"b69" => data <= x"2c";
            when "00" & x"b6a" => data <= x"e6";
            when "00" & x"b6b" => data <= x"fe";
            when "00" & x"b6c" => data <= x"50";
            when "00" & x"b6d" => data <= x"fb";
            when "00" & x"b6e" => data <= x"b0";
            when "00" & x"b6f" => data <= x"0d";
            when "00" & x"b70" => data <= x"e0";
            when "00" & x"b71" => data <= x"04";
            when "00" & x"b72" => data <= x"d0";
            when "00" & x"b73" => data <= x"11";
            when "00" & x"b74" => data <= x"20";
            when "00" & x"b75" => data <= x"14";
            when "00" & x"b76" => data <= x"04";
            when "00" & x"b77" => data <= x"20";
            when "00" & x"b78" => data <= x"95";
            when "00" & x"b79" => data <= x"06";
            when "00" & x"b7a" => data <= x"4c";
            when "00" & x"b7b" => data <= x"32";
            when "00" & x"b7c" => data <= x"00";
            when "00" & x"b7d" => data <= x"4a";
            when "00" & x"b7e" => data <= x"90";
            when "00" & x"b7f" => data <= x"05";
            when "00" & x"b80" => data <= x"a0";
            when "00" & x"b81" => data <= x"88";
            when "00" & x"b82" => data <= x"8c";
            when "00" & x"b83" => data <= x"e0";
            when "00" & x"b84" => data <= x"fe";
            when "00" & x"b85" => data <= x"28";
            when "00" & x"b86" => data <= x"60";
            when "00" & x"b87" => data <= x"58";
            when "00" & x"b88" => data <= x"b0";
            when "00" & x"b89" => data <= x"11";
            when "00" & x"b8a" => data <= x"d0";
            when "00" & x"b8b" => data <= x"03";
            when "00" & x"b8c" => data <= x"4c";
            when "00" & x"b8d" => data <= x"9c";
            when "00" & x"b8e" => data <= x"05";
            when "00" & x"b8f" => data <= x"a2";
            when "00" & x"b90" => data <= x"00";
            when "00" & x"b91" => data <= x"a0";
            when "00" & x"b92" => data <= x"ff";
            when "00" & x"b93" => data <= x"a9";
            when "00" & x"b94" => data <= x"fd";
            when "00" & x"b95" => data <= x"20";
            when "00" & x"b96" => data <= x"f4";
            when "00" & x"b97" => data <= x"ff";
            when "00" & x"b98" => data <= x"8a";
            when "00" & x"b99" => data <= x"f0";
            when "00" & x"b9a" => data <= x"d9";
            when "00" & x"b9b" => data <= x"a9";
            when "00" & x"b9c" => data <= x"ff";
            when "00" & x"b9d" => data <= x"20";
            when "00" & x"b9e" => data <= x"06";
            when "00" & x"b9f" => data <= x"04";
            when "00" & x"ba0" => data <= x"90";
            when "00" & x"ba1" => data <= x"f9";
            when "00" & x"ba2" => data <= x"20";
            when "00" & x"ba3" => data <= x"d2";
            when "00" & x"ba4" => data <= x"04";
            when "00" & x"ba5" => data <= x"a9";
            when "00" & x"ba6" => data <= x"07";
            when "00" & x"ba7" => data <= x"20";
            when "00" & x"ba8" => data <= x"cb";
            when "00" & x"ba9" => data <= x"04";
            when "00" & x"baa" => data <= x"a0";
            when "00" & x"bab" => data <= x"00";
            when "00" & x"bac" => data <= x"84";
            when "00" & x"bad" => data <= x"00";
            when "00" & x"bae" => data <= x"b1";
            when "00" & x"baf" => data <= x"00";
            when "00" & x"bb0" => data <= x"8d";
            when "00" & x"bb1" => data <= x"e5";
            when "00" & x"bb2" => data <= x"fe";
            when "00" & x"bb3" => data <= x"ea";
            when "00" & x"bb4" => data <= x"ea";
            when "00" & x"bb5" => data <= x"ea";
            when "00" & x"bb6" => data <= x"c8";
            when "00" & x"bb7" => data <= x"d0";
            when "00" & x"bb8" => data <= x"f5";
            when "00" & x"bb9" => data <= x"e6";
            when "00" & x"bba" => data <= x"54";
            when "00" & x"bbb" => data <= x"d0";
            when "00" & x"bbc" => data <= x"06";
            when "00" & x"bbd" => data <= x"e6";
            when "00" & x"bbe" => data <= x"55";
            when "00" & x"bbf" => data <= x"d0";
            when "00" & x"bc0" => data <= x"02";
            when "00" & x"bc1" => data <= x"e6";
            when "00" & x"bc2" => data <= x"56";
            when "00" & x"bc3" => data <= x"e6";
            when "00" & x"bc4" => data <= x"01";
            when "00" & x"bc5" => data <= x"24";
            when "00" & x"bc6" => data <= x"01";
            when "00" & x"bc7" => data <= x"50";
            when "00" & x"bc8" => data <= x"dc";
            when "00" & x"bc9" => data <= x"20";
            when "00" & x"bca" => data <= x"d2";
            when "00" & x"bcb" => data <= x"04";
            when "00" & x"bcc" => data <= x"a9";
            when "00" & x"bcd" => data <= x"04";
            when "00" & x"bce" => data <= x"a0";
            when "00" & x"bcf" => data <= x"00";
            when "00" & x"bd0" => data <= x"a2";
            when "00" & x"bd1" => data <= x"53";
            when "00" & x"bd2" => data <= x"4c";
            when "00" & x"bd3" => data <= x"06";
            when "00" & x"bd4" => data <= x"04";
            when "00" & x"bd5" => data <= x"a9";
            when "00" & x"bd6" => data <= x"80";
            when "00" & x"bd7" => data <= x"85";
            when "00" & x"bd8" => data <= x"54";
            when "00" & x"bd9" => data <= x"85";
            when "00" & x"bda" => data <= x"01";
            when "00" & x"bdb" => data <= x"a9";
            when "00" & x"bdc" => data <= x"20";
            when "00" & x"bdd" => data <= x"2d";
            when "00" & x"bde" => data <= x"06";
            when "00" & x"bdf" => data <= x"80";
            when "00" & x"be0" => data <= x"a8";
            when "00" & x"be1" => data <= x"84";
            when "00" & x"be2" => data <= x"53";
            when "00" & x"be3" => data <= x"f0";
            when "00" & x"be4" => data <= x"19";
            when "00" & x"be5" => data <= x"ae";
            when "00" & x"be6" => data <= x"07";
            when "00" & x"be7" => data <= x"80";
            when "00" & x"be8" => data <= x"e8";
            when "00" & x"be9" => data <= x"bd";
            when "00" & x"bea" => data <= x"00";
            when "00" & x"beb" => data <= x"80";
            when "00" & x"bec" => data <= x"d0";
            when "00" & x"bed" => data <= x"fa";
            when "00" & x"bee" => data <= x"bd";
            when "00" & x"bef" => data <= x"01";
            when "00" & x"bf0" => data <= x"80";
            when "00" & x"bf1" => data <= x"85";
            when "00" & x"bf2" => data <= x"53";
            when "00" & x"bf3" => data <= x"bd";
            when "00" & x"bf4" => data <= x"02";
            when "00" & x"bf5" => data <= x"80";
            when "00" & x"bf6" => data <= x"85";
            when "00" & x"bf7" => data <= x"54";
            when "00" & x"bf8" => data <= x"bc";
            when "00" & x"bf9" => data <= x"03";
            when "00" & x"bfa" => data <= x"80";
            when "00" & x"bfb" => data <= x"bd";
            when "00" & x"bfc" => data <= x"04";
            when "00" & x"bfd" => data <= x"80";
            when "00" & x"bfe" => data <= x"85";
            when "00" & x"bff" => data <= x"56";
            when "00" & x"c00" => data <= x"84";
            when "00" & x"c01" => data <= x"55";
            when "00" & x"c02" => data <= x"60";
            when "00" & x"c03" => data <= x"37";
            when "00" & x"c04" => data <= x"05";
            when "00" & x"c05" => data <= x"96";
            when "00" & x"c06" => data <= x"05";
            when "00" & x"c07" => data <= x"f2";
            when "00" & x"c08" => data <= x"05";
            when "00" & x"c09" => data <= x"07";
            when "00" & x"c0a" => data <= x"06";
            when "00" & x"c0b" => data <= x"27";
            when "00" & x"c0c" => data <= x"06";
            when "00" & x"c0d" => data <= x"68";
            when "00" & x"c0e" => data <= x"06";
            when "00" & x"c0f" => data <= x"5e";
            when "00" & x"c10" => data <= x"05";
            when "00" & x"c11" => data <= x"2d";
            when "00" & x"c12" => data <= x"05";
            when "00" & x"c13" => data <= x"20";
            when "00" & x"c14" => data <= x"05";
            when "00" & x"c15" => data <= x"42";
            when "00" & x"c16" => data <= x"05";
            when "00" & x"c17" => data <= x"a9";
            when "00" & x"c18" => data <= x"05";
            when "00" & x"c19" => data <= x"d1";
            when "00" & x"c1a" => data <= x"05";
            when "00" & x"c1b" => data <= x"86";
            when "00" & x"c1c" => data <= x"88";
            when "00" & x"c1d" => data <= x"96";
            when "00" & x"c1e" => data <= x"98";
            when "00" & x"c1f" => data <= x"18";
            when "00" & x"c20" => data <= x"18";
            when "00" & x"c21" => data <= x"82";
            when "00" & x"c22" => data <= x"18";
            when "00" & x"c23" => data <= x"20";
            when "00" & x"c24" => data <= x"c5";
            when "00" & x"c25" => data <= x"06";
            when "00" & x"c26" => data <= x"a8";
            when "00" & x"c27" => data <= x"20";
            when "00" & x"c28" => data <= x"c5";
            when "00" & x"c29" => data <= x"06";
            when "00" & x"c2a" => data <= x"20";
            when "00" & x"c2b" => data <= x"d4";
            when "00" & x"c2c" => data <= x"ff";
            when "00" & x"c2d" => data <= x"4c";
            when "00" & x"c2e" => data <= x"9c";
            when "00" & x"c2f" => data <= x"05";
            when "00" & x"c30" => data <= x"20";
            when "00" & x"c31" => data <= x"c5";
            when "00" & x"c32" => data <= x"06";
            when "00" & x"c33" => data <= x"a8";
            when "00" & x"c34" => data <= x"20";
            when "00" & x"c35" => data <= x"d7";
            when "00" & x"c36" => data <= x"ff";
            when "00" & x"c37" => data <= x"4c";
            when "00" & x"c38" => data <= x"3a";
            when "00" & x"c39" => data <= x"05";
            when "00" & x"c3a" => data <= x"20";
            when "00" & x"c3b" => data <= x"e0";
            when "00" & x"c3c" => data <= x"ff";
            when "00" & x"c3d" => data <= x"6a";
            when "00" & x"c3e" => data <= x"20";
            when "00" & x"c3f" => data <= x"95";
            when "00" & x"c40" => data <= x"06";
            when "00" & x"c41" => data <= x"2a";
            when "00" & x"c42" => data <= x"4c";
            when "00" & x"c43" => data <= x"9e";
            when "00" & x"c44" => data <= x"05";
            when "00" & x"c45" => data <= x"20";
            when "00" & x"c46" => data <= x"c5";
            when "00" & x"c47" => data <= x"06";
            when "00" & x"c48" => data <= x"f0";
            when "00" & x"c49" => data <= x"0b";
            when "00" & x"c4a" => data <= x"48";
            when "00" & x"c4b" => data <= x"20";
            when "00" & x"c4c" => data <= x"82";
            when "00" & x"c4d" => data <= x"05";
            when "00" & x"c4e" => data <= x"68";
            when "00" & x"c4f" => data <= x"20";
            when "00" & x"c50" => data <= x"ce";
            when "00" & x"c51" => data <= x"ff";
            when "00" & x"c52" => data <= x"4c";
            when "00" & x"c53" => data <= x"9e";
            when "00" & x"c54" => data <= x"05";
            when "00" & x"c55" => data <= x"20";
            when "00" & x"c56" => data <= x"c5";
            when "00" & x"c57" => data <= x"06";
            when "00" & x"c58" => data <= x"a8";
            when "00" & x"c59" => data <= x"a9";
            when "00" & x"c5a" => data <= x"00";
            when "00" & x"c5b" => data <= x"20";
            when "00" & x"c5c" => data <= x"ce";
            when "00" & x"c5d" => data <= x"ff";
            when "00" & x"c5e" => data <= x"4c";
            when "00" & x"c5f" => data <= x"9c";
            when "00" & x"c60" => data <= x"05";
            when "00" & x"c61" => data <= x"20";
            when "00" & x"c62" => data <= x"c5";
            when "00" & x"c63" => data <= x"06";
            when "00" & x"c64" => data <= x"a8";
            when "00" & x"c65" => data <= x"a2";
            when "00" & x"c66" => data <= x"04";
            when "00" & x"c67" => data <= x"20";
            when "00" & x"c68" => data <= x"c5";
            when "00" & x"c69" => data <= x"06";
            when "00" & x"c6a" => data <= x"95";
            when "00" & x"c6b" => data <= x"ff";
            when "00" & x"c6c" => data <= x"ca";
            when "00" & x"c6d" => data <= x"d0";
            when "00" & x"c6e" => data <= x"f8";
            when "00" & x"c6f" => data <= x"20";
            when "00" & x"c70" => data <= x"c5";
            when "00" & x"c71" => data <= x"06";
            when "00" & x"c72" => data <= x"20";
            when "00" & x"c73" => data <= x"da";
            when "00" & x"c74" => data <= x"ff";
            when "00" & x"c75" => data <= x"20";
            when "00" & x"c76" => data <= x"95";
            when "00" & x"c77" => data <= x"06";
            when "00" & x"c78" => data <= x"a2";
            when "00" & x"c79" => data <= x"03";
            when "00" & x"c7a" => data <= x"b5";
            when "00" & x"c7b" => data <= x"00";
            when "00" & x"c7c" => data <= x"20";
            when "00" & x"c7d" => data <= x"95";
            when "00" & x"c7e" => data <= x"06";
            when "00" & x"c7f" => data <= x"ca";
            when "00" & x"c80" => data <= x"10";
            when "00" & x"c81" => data <= x"f8";
            when "00" & x"c82" => data <= x"4c";
            when "00" & x"c83" => data <= x"36";
            when "00" & x"c84" => data <= x"00";
            when "00" & x"c85" => data <= x"a2";
            when "00" & x"c86" => data <= x"00";
            when "00" & x"c87" => data <= x"a0";
            when "00" & x"c88" => data <= x"00";
            when "00" & x"c89" => data <= x"20";
            when "00" & x"c8a" => data <= x"c5";
            when "00" & x"c8b" => data <= x"06";
            when "00" & x"c8c" => data <= x"99";
            when "00" & x"c8d" => data <= x"00";
            when "00" & x"c8e" => data <= x"07";
            when "00" & x"c8f" => data <= x"c8";
            when "00" & x"c90" => data <= x"f0";
            when "00" & x"c91" => data <= x"04";
            when "00" & x"c92" => data <= x"c9";
            when "00" & x"c93" => data <= x"0d";
            when "00" & x"c94" => data <= x"d0";
            when "00" & x"c95" => data <= x"f3";
            when "00" & x"c96" => data <= x"a0";
            when "00" & x"c97" => data <= x"07";
            when "00" & x"c98" => data <= x"60";
            when "00" & x"c99" => data <= x"20";
            when "00" & x"c9a" => data <= x"82";
            when "00" & x"c9b" => data <= x"05";
            when "00" & x"c9c" => data <= x"20";
            when "00" & x"c9d" => data <= x"f7";
            when "00" & x"c9e" => data <= x"ff";
            when "00" & x"c9f" => data <= x"a9";
            when "00" & x"ca0" => data <= x"7f";
            when "00" & x"ca1" => data <= x"2c";
            when "00" & x"ca2" => data <= x"e2";
            when "00" & x"ca3" => data <= x"fe";
            when "00" & x"ca4" => data <= x"50";
            when "00" & x"ca5" => data <= x"fb";
            when "00" & x"ca6" => data <= x"8d";
            when "00" & x"ca7" => data <= x"e3";
            when "00" & x"ca8" => data <= x"fe";
            when "00" & x"ca9" => data <= x"4c";
            when "00" & x"caa" => data <= x"36";
            when "00" & x"cab" => data <= x"00";
            when "00" & x"cac" => data <= x"a2";
            when "00" & x"cad" => data <= x"10";
            when "00" & x"cae" => data <= x"20";
            when "00" & x"caf" => data <= x"c5";
            when "00" & x"cb0" => data <= x"06";
            when "00" & x"cb1" => data <= x"95";
            when "00" & x"cb2" => data <= x"01";
            when "00" & x"cb3" => data <= x"ca";
            when "00" & x"cb4" => data <= x"d0";
            when "00" & x"cb5" => data <= x"f8";
            when "00" & x"cb6" => data <= x"20";
            when "00" & x"cb7" => data <= x"82";
            when "00" & x"cb8" => data <= x"05";
            when "00" & x"cb9" => data <= x"86";
            when "00" & x"cba" => data <= x"00";
            when "00" & x"cbb" => data <= x"84";
            when "00" & x"cbc" => data <= x"01";
            when "00" & x"cbd" => data <= x"a0";
            when "00" & x"cbe" => data <= x"00";
            when "00" & x"cbf" => data <= x"20";
            when "00" & x"cc0" => data <= x"c5";
            when "00" & x"cc1" => data <= x"06";
            when "00" & x"cc2" => data <= x"20";
            when "00" & x"cc3" => data <= x"dd";
            when "00" & x"cc4" => data <= x"ff";
            when "00" & x"cc5" => data <= x"20";
            when "00" & x"cc6" => data <= x"95";
            when "00" & x"cc7" => data <= x"06";
            when "00" & x"cc8" => data <= x"a2";
            when "00" & x"cc9" => data <= x"10";
            when "00" & x"cca" => data <= x"b5";
            when "00" & x"ccb" => data <= x"01";
            when "00" & x"ccc" => data <= x"20";
            when "00" & x"ccd" => data <= x"95";
            when "00" & x"cce" => data <= x"06";
            when "00" & x"ccf" => data <= x"ca";
            when "00" & x"cd0" => data <= x"d0";
            when "00" & x"cd1" => data <= x"f8";
            when "00" & x"cd2" => data <= x"f0";
            when "00" & x"cd3" => data <= x"d5";
            when "00" & x"cd4" => data <= x"a2";
            when "00" & x"cd5" => data <= x"0d";
            when "00" & x"cd6" => data <= x"20";
            when "00" & x"cd7" => data <= x"c5";
            when "00" & x"cd8" => data <= x"06";
            when "00" & x"cd9" => data <= x"95";
            when "00" & x"cda" => data <= x"ff";
            when "00" & x"cdb" => data <= x"ca";
            when "00" & x"cdc" => data <= x"d0";
            when "00" & x"cdd" => data <= x"f8";
            when "00" & x"cde" => data <= x"20";
            when "00" & x"cdf" => data <= x"c5";
            when "00" & x"ce0" => data <= x"06";
            when "00" & x"ce1" => data <= x"a0";
            when "00" & x"ce2" => data <= x"00";
            when "00" & x"ce3" => data <= x"20";
            when "00" & x"ce4" => data <= x"d1";
            when "00" & x"ce5" => data <= x"ff";
            when "00" & x"ce6" => data <= x"48";
            when "00" & x"ce7" => data <= x"a2";
            when "00" & x"ce8" => data <= x"0c";
            when "00" & x"ce9" => data <= x"b5";
            when "00" & x"cea" => data <= x"00";
            when "00" & x"ceb" => data <= x"20";
            when "00" & x"cec" => data <= x"95";
            when "00" & x"ced" => data <= x"06";
            when "00" & x"cee" => data <= x"ca";
            when "00" & x"cef" => data <= x"10";
            when "00" & x"cf0" => data <= x"f8";
            when "00" & x"cf1" => data <= x"68";
            when "00" & x"cf2" => data <= x"4c";
            when "00" & x"cf3" => data <= x"3a";
            when "00" & x"cf4" => data <= x"05";
            when "00" & x"cf5" => data <= x"20";
            when "00" & x"cf6" => data <= x"c5";
            when "00" & x"cf7" => data <= x"06";
            when "00" & x"cf8" => data <= x"aa";
            when "00" & x"cf9" => data <= x"20";
            when "00" & x"cfa" => data <= x"c5";
            when "00" & x"cfb" => data <= x"06";
            when "00" & x"cfc" => data <= x"20";
            when "00" & x"cfd" => data <= x"f4";
            when "00" & x"cfe" => data <= x"ff";
            when "00" & x"cff" => data <= x"2c";
            when "00" & x"d00" => data <= x"e2";
            when "00" & x"d01" => data <= x"fe";
            when "00" & x"d02" => data <= x"50";
            when "00" & x"d03" => data <= x"fb";
            when "00" & x"d04" => data <= x"8e";
            when "00" & x"d05" => data <= x"e3";
            when "00" & x"d06" => data <= x"fe";
            when "00" & x"d07" => data <= x"4c";
            when "00" & x"d08" => data <= x"36";
            when "00" & x"d09" => data <= x"00";
            when "00" & x"d0a" => data <= x"20";
            when "00" & x"d0b" => data <= x"c5";
            when "00" & x"d0c" => data <= x"06";
            when "00" & x"d0d" => data <= x"aa";
            when "00" & x"d0e" => data <= x"20";
            when "00" & x"d0f" => data <= x"c5";
            when "00" & x"d10" => data <= x"06";
            when "00" & x"d11" => data <= x"a8";
            when "00" & x"d12" => data <= x"20";
            when "00" & x"d13" => data <= x"c5";
            when "00" & x"d14" => data <= x"06";
            when "00" & x"d15" => data <= x"20";
            when "00" & x"d16" => data <= x"f4";
            when "00" & x"d17" => data <= x"ff";
            when "00" & x"d18" => data <= x"49";
            when "00" & x"d19" => data <= x"9d";
            when "00" & x"d1a" => data <= x"f0";
            when "00" & x"d1b" => data <= x"eb";
            when "00" & x"d1c" => data <= x"6a";
            when "00" & x"d1d" => data <= x"20";
            when "00" & x"d1e" => data <= x"95";
            when "00" & x"d1f" => data <= x"06";
            when "00" & x"d20" => data <= x"2c";
            when "00" & x"d21" => data <= x"e2";
            when "00" & x"d22" => data <= x"fe";
            when "00" & x"d23" => data <= x"50";
            when "00" & x"d24" => data <= x"fb";
            when "00" & x"d25" => data <= x"8c";
            when "00" & x"d26" => data <= x"e3";
            when "00" & x"d27" => data <= x"fe";
            when "00" & x"d28" => data <= x"70";
            when "00" & x"d29" => data <= x"d5";
            when "00" & x"d2a" => data <= x"20";
            when "00" & x"d2b" => data <= x"c5";
            when "00" & x"d2c" => data <= x"06";
            when "00" & x"d2d" => data <= x"a8";
            when "00" & x"d2e" => data <= x"2c";
            when "00" & x"d2f" => data <= x"e2";
            when "00" & x"d30" => data <= x"fe";
            when "00" & x"d31" => data <= x"10";
            when "00" & x"d32" => data <= x"fb";
            when "00" & x"d33" => data <= x"ae";
            when "00" & x"d34" => data <= x"e3";
            when "00" & x"d35" => data <= x"fe";
            when "00" & x"d36" => data <= x"ca";
            when "00" & x"d37" => data <= x"30";
            when "00" & x"d38" => data <= x"0f";
            when "00" & x"d39" => data <= x"2c";
            when "00" & x"d3a" => data <= x"e2";
            when "00" & x"d3b" => data <= x"fe";
            when "00" & x"d3c" => data <= x"10";
            when "00" & x"d3d" => data <= x"fb";
            when "00" & x"d3e" => data <= x"ad";
            when "00" & x"d3f" => data <= x"e3";
            when "00" & x"d40" => data <= x"fe";
            when "00" & x"d41" => data <= x"9d";
            when "00" & x"d42" => data <= x"28";
            when "00" & x"d43" => data <= x"01";
            when "00" & x"d44" => data <= x"ca";
            when "00" & x"d45" => data <= x"10";
            when "00" & x"d46" => data <= x"f2";
            when "00" & x"d47" => data <= x"98";
            when "00" & x"d48" => data <= x"a2";
            when "00" & x"d49" => data <= x"28";
            when "00" & x"d4a" => data <= x"a0";
            when "00" & x"d4b" => data <= x"01";
            when "00" & x"d4c" => data <= x"20";
            when "00" & x"d4d" => data <= x"f1";
            when "00" & x"d4e" => data <= x"ff";
            when "00" & x"d4f" => data <= x"2c";
            when "00" & x"d50" => data <= x"e2";
            when "00" & x"d51" => data <= x"fe";
            when "00" & x"d52" => data <= x"10";
            when "00" & x"d53" => data <= x"fb";
            when "00" & x"d54" => data <= x"ae";
            when "00" & x"d55" => data <= x"e3";
            when "00" & x"d56" => data <= x"fe";
            when "00" & x"d57" => data <= x"ca";
            when "00" & x"d58" => data <= x"30";
            when "00" & x"d59" => data <= x"0e";
            when "00" & x"d5a" => data <= x"bc";
            when "00" & x"d5b" => data <= x"28";
            when "00" & x"d5c" => data <= x"01";
            when "00" & x"d5d" => data <= x"2c";
            when "00" & x"d5e" => data <= x"e2";
            when "00" & x"d5f" => data <= x"fe";
            when "00" & x"d60" => data <= x"50";
            when "00" & x"d61" => data <= x"fb";
            when "00" & x"d62" => data <= x"8c";
            when "00" & x"d63" => data <= x"e3";
            when "00" & x"d64" => data <= x"fe";
            when "00" & x"d65" => data <= x"ca";
            when "00" & x"d66" => data <= x"10";
            when "00" & x"d67" => data <= x"f2";
            when "00" & x"d68" => data <= x"4c";
            when "00" & x"d69" => data <= x"36";
            when "00" & x"d6a" => data <= x"00";
            when "00" & x"d6b" => data <= x"a2";
            when "00" & x"d6c" => data <= x"04";
            when "00" & x"d6d" => data <= x"20";
            when "00" & x"d6e" => data <= x"c5";
            when "00" & x"d6f" => data <= x"06";
            when "00" & x"d70" => data <= x"95";
            when "00" & x"d71" => data <= x"00";
            when "00" & x"d72" => data <= x"ca";
            when "00" & x"d73" => data <= x"10";
            when "00" & x"d74" => data <= x"f8";
            when "00" & x"d75" => data <= x"e8";
            when "00" & x"d76" => data <= x"a0";
            when "00" & x"d77" => data <= x"00";
            when "00" & x"d78" => data <= x"8a";
            when "00" & x"d79" => data <= x"20";
            when "00" & x"d7a" => data <= x"f1";
            when "00" & x"d7b" => data <= x"ff";
            when "00" & x"d7c" => data <= x"90";
            when "00" & x"d7d" => data <= x"05";
            when "00" & x"d7e" => data <= x"a9";
            when "00" & x"d7f" => data <= x"ff";
            when "00" & x"d80" => data <= x"4c";
            when "00" & x"d81" => data <= x"9e";
            when "00" & x"d82" => data <= x"05";
            when "00" & x"d83" => data <= x"a2";
            when "00" & x"d84" => data <= x"00";
            when "00" & x"d85" => data <= x"a9";
            when "00" & x"d86" => data <= x"7f";
            when "00" & x"d87" => data <= x"20";
            when "00" & x"d88" => data <= x"95";
            when "00" & x"d89" => data <= x"06";
            when "00" & x"d8a" => data <= x"bd";
            when "00" & x"d8b" => data <= x"00";
            when "00" & x"d8c" => data <= x"07";
            when "00" & x"d8d" => data <= x"20";
            when "00" & x"d8e" => data <= x"95";
            when "00" & x"d8f" => data <= x"06";
            when "00" & x"d90" => data <= x"e8";
            when "00" & x"d91" => data <= x"c9";
            when "00" & x"d92" => data <= x"0d";
            when "00" & x"d93" => data <= x"d0";
            when "00" & x"d94" => data <= x"f5";
            when "00" & x"d95" => data <= x"4c";
            when "00" & x"d96" => data <= x"36";
            when "00" & x"d97" => data <= x"00";
            when "00" & x"d98" => data <= x"2c";
            when "00" & x"d99" => data <= x"e2";
            when "00" & x"d9a" => data <= x"fe";
            when "00" & x"d9b" => data <= x"50";
            when "00" & x"d9c" => data <= x"fb";
            when "00" & x"d9d" => data <= x"8d";
            when "00" & x"d9e" => data <= x"e3";
            when "00" & x"d9f" => data <= x"fe";
            when "00" & x"da0" => data <= x"60";
            when "00" & x"da1" => data <= x"2c";
            when "00" & x"da2" => data <= x"e6";
            when "00" & x"da3" => data <= x"fe";
            when "00" & x"da4" => data <= x"50";
            when "00" & x"da5" => data <= x"fb";
            when "00" & x"da6" => data <= x"8d";
            when "00" & x"da7" => data <= x"e7";
            when "00" & x"da8" => data <= x"fe";
            when "00" & x"da9" => data <= x"60";
            when "00" & x"daa" => data <= x"a5";
            when "00" & x"dab" => data <= x"ff";
            when "00" & x"dac" => data <= x"38";
            when "00" & x"dad" => data <= x"6a";
            when "00" & x"dae" => data <= x"30";
            when "00" & x"daf" => data <= x"0f";
            when "00" & x"db0" => data <= x"48";
            when "00" & x"db1" => data <= x"a9";
            when "00" & x"db2" => data <= x"00";
            when "00" & x"db3" => data <= x"20";
            when "00" & x"db4" => data <= x"bc";
            when "00" & x"db5" => data <= x"06";
            when "00" & x"db6" => data <= x"98";
            when "00" & x"db7" => data <= x"20";
            when "00" & x"db8" => data <= x"bc";
            when "00" & x"db9" => data <= x"06";
            when "00" & x"dba" => data <= x"8a";
            when "00" & x"dbb" => data <= x"20";
            when "00" & x"dbc" => data <= x"bc";
            when "00" & x"dbd" => data <= x"06";
            when "00" & x"dbe" => data <= x"68";
            when "00" & x"dbf" => data <= x"2c";
            when "00" & x"dc0" => data <= x"e0";
            when "00" & x"dc1" => data <= x"fe";
            when "00" & x"dc2" => data <= x"50";
            when "00" & x"dc3" => data <= x"fb";
            when "00" & x"dc4" => data <= x"8d";
            when "00" & x"dc5" => data <= x"e1";
            when "00" & x"dc6" => data <= x"fe";
            when "00" & x"dc7" => data <= x"60";
            when "00" & x"dc8" => data <= x"2c";
            when "00" & x"dc9" => data <= x"e2";
            when "00" & x"dca" => data <= x"fe";
            when "00" & x"dcb" => data <= x"10";
            when "00" & x"dcc" => data <= x"fb";
            when "00" & x"dcd" => data <= x"ad";
            when "00" & x"dce" => data <= x"e3";
            when "00" & x"dcf" => data <= x"fe";
            when "00" & x"dd0" => data <= x"60";
            when "00" & x"dd1" => data <= x"00";
            when "00" & x"dd2" => data <= x"00";
            when "00" & x"dd3" => data <= x"00";
            when "00" & x"dd4" => data <= x"00";
            when "00" & x"dd5" => data <= x"00";
            when "00" & x"dd6" => data <= x"00";
            when "00" & x"dd7" => data <= x"00";
            when "00" & x"dd8" => data <= x"00";
            when "00" & x"dd9" => data <= x"00";
            when "00" & x"dda" => data <= x"00";
            when "00" & x"ddb" => data <= x"00";
            when "00" & x"ddc" => data <= x"00";
            when "00" & x"ddd" => data <= x"a2";
            when "00" & x"dde" => data <= x"11";
            when "00" & x"ddf" => data <= x"a0";
            when "00" & x"de0" => data <= x"13";
            when "00" & x"de1" => data <= x"60";
            when "00" & x"de2" => data <= x"20";
            when "00" & x"de3" => data <= x"e1";
            when "00" & x"de4" => data <= x"83";
            when "00" & x"de5" => data <= x"a9";
            when "00" & x"de6" => data <= x"77";
            when "00" & x"de7" => data <= x"4c";
            when "00" & x"de8" => data <= x"f4";
            when "00" & x"de9" => data <= x"ff";
            when "00" & x"dea" => data <= x"20";
            when "00" & x"deb" => data <= x"e2";
            when "00" & x"dec" => data <= x"8d";
            when "00" & x"ded" => data <= x"a9";
            when "00" & x"dee" => data <= x"00";
            when "00" & x"def" => data <= x"18";
            when "00" & x"df0" => data <= x"69";
            when "00" & x"df1" => data <= x"20";
            when "00" & x"df2" => data <= x"f0";
            when "00" & x"df3" => data <= x"ed";
            when "00" & x"df4" => data <= x"a8";
            when "00" & x"df5" => data <= x"20";
            when "00" & x"df6" => data <= x"05";
            when "00" & x"df7" => data <= x"8e";
            when "00" & x"df8" => data <= x"d0";
            when "00" & x"df9" => data <= x"f5";
            when "00" & x"dfa" => data <= x"98";
            when "00" & x"dfb" => data <= x"f0";
            when "00" & x"dfc" => data <= x"ed";
            when "00" & x"dfd" => data <= x"20";
            when "00" & x"dfe" => data <= x"7b";
            when "00" & x"dff" => data <= x"90";
            when "00" & x"e00" => data <= x"90";
            when "00" & x"e01" => data <= x"03";
            when "00" & x"e02" => data <= x"4c";
            when "00" & x"e03" => data <= x"ad";
            when "00" & x"e04" => data <= x"90";
            when "00" & x"e05" => data <= x"48";
            when "00" & x"e06" => data <= x"20";
            when "00" & x"e07" => data <= x"51";
            when "00" & x"e08" => data <= x"90";
            when "00" & x"e09" => data <= x"b0";
            when "00" & x"e0a" => data <= x"45";
            when "00" & x"e0b" => data <= x"b9";
            when "00" & x"e0c" => data <= x"1b";
            when "00" & x"e0d" => data <= x"11";
            when "00" & x"e0e" => data <= x"49";
            when "00" & x"e0f" => data <= x"ff";
            when "00" & x"e10" => data <= x"2d";
            when "00" & x"e11" => data <= x"c0";
            when "00" & x"e12" => data <= x"10";
            when "00" & x"e13" => data <= x"8d";
            when "00" & x"e14" => data <= x"c0";
            when "00" & x"e15" => data <= x"10";
            when "00" & x"e16" => data <= x"b9";
            when "00" & x"e17" => data <= x"17";
            when "00" & x"e18" => data <= x"11";
            when "00" & x"e19" => data <= x"29";
            when "00" & x"e1a" => data <= x"60";
            when "00" & x"e1b" => data <= x"f0";
            when "00" & x"e1c" => data <= x"33";
            when "00" & x"e1d" => data <= x"20";
            when "00" & x"e1e" => data <= x"55";
            when "00" & x"e1f" => data <= x"8e";
            when "00" & x"e20" => data <= x"b9";
            when "00" & x"e21" => data <= x"17";
            when "00" & x"e22" => data <= x"11";
            when "00" & x"e23" => data <= x"29";
            when "00" & x"e24" => data <= x"20";
            when "00" & x"e25" => data <= x"f0";
            when "00" & x"e26" => data <= x"26";
            when "00" & x"e27" => data <= x"ae";
            when "00" & x"e28" => data <= x"c4";
            when "00" & x"e29" => data <= x"10";
            when "00" & x"e2a" => data <= x"b9";
            when "00" & x"e2b" => data <= x"14";
            when "00" & x"e2c" => data <= x"11";
            when "00" & x"e2d" => data <= x"9d";
            when "00" & x"e2e" => data <= x"0c";
            when "00" & x"e2f" => data <= x"0f";
            when "00" & x"e30" => data <= x"b9";
            when "00" & x"e31" => data <= x"15";
            when "00" & x"e32" => data <= x"11";
            when "00" & x"e33" => data <= x"9d";
            when "00" & x"e34" => data <= x"0d";
            when "00" & x"e35" => data <= x"0f";
            when "00" & x"e36" => data <= x"b9";
            when "00" & x"e37" => data <= x"16";
            when "00" & x"e38" => data <= x"11";
            when "00" & x"e39" => data <= x"20";
            when "00" & x"e3a" => data <= x"0b";
            when "00" & x"e3b" => data <= x"82";
            when "00" & x"e3c" => data <= x"5d";
            when "00" & x"e3d" => data <= x"0e";
            when "00" & x"e3e" => data <= x"0f";
            when "00" & x"e3f" => data <= x"29";
            when "00" & x"e40" => data <= x"30";
            when "00" & x"e41" => data <= x"5d";
            when "00" & x"e42" => data <= x"0e";
            when "00" & x"e43" => data <= x"0f";
            when "00" & x"e44" => data <= x"9d";
            when "00" & x"e45" => data <= x"0e";
            when "00" & x"e46" => data <= x"0f";
            when "00" & x"e47" => data <= x"20";
            when "00" & x"e48" => data <= x"b4";
            when "00" & x"e49" => data <= x"8a";
            when "00" & x"e4a" => data <= x"ac";
            when "00" & x"e4b" => data <= x"c2";
            when "00" & x"e4c" => data <= x"10";
            when "00" & x"e4d" => data <= x"20";
            when "00" & x"e4e" => data <= x"4b";
            when "00" & x"e4f" => data <= x"91";
            when "00" & x"e50" => data <= x"ae";
            when "00" & x"e51" => data <= x"c6";
            when "00" & x"e52" => data <= x"10";
            when "00" & x"e53" => data <= x"68";
            when "00" & x"e54" => data <= x"60";
            when "00" & x"e55" => data <= x"20";
            when "00" & x"e56" => data <= x"83";
            when "00" & x"e57" => data <= x"8e";
            when "00" & x"e58" => data <= x"a2";
            when "00" & x"e59" => data <= x"07";
            when "00" & x"e5a" => data <= x"b9";
            when "00" & x"e5b" => data <= x"0c";
            when "00" & x"e5c" => data <= x"11";
            when "00" & x"e5d" => data <= x"95";
            when "00" & x"e5e" => data <= x"c6";
            when "00" & x"e5f" => data <= x"88";
            when "00" & x"e60" => data <= x"88";
            when "00" & x"e61" => data <= x"ca";
            when "00" & x"e62" => data <= x"d0";
            when "00" & x"e63" => data <= x"f6";
            when "00" & x"e64" => data <= x"20";
            when "00" & x"e65" => data <= x"96";
            when "00" & x"e66" => data <= x"82";
            when "00" & x"e67" => data <= x"90";
            when "00" & x"e68" => data <= x"27";
            when "00" & x"e69" => data <= x"8c";
            when "00" & x"e6a" => data <= x"c4";
            when "00" & x"e6b" => data <= x"10";
            when "00" & x"e6c" => data <= x"b9";
            when "00" & x"e6d" => data <= x"0e";
            when "00" & x"e6e" => data <= x"0f";
            when "00" & x"e6f" => data <= x"be";
            when "00" & x"e70" => data <= x"0f";
            when "00" & x"e71" => data <= x"0f";
            when "00" & x"e72" => data <= x"ac";
            when "00" & x"e73" => data <= x"c2";
            when "00" & x"e74" => data <= x"10";
            when "00" & x"e75" => data <= x"59";
            when "00" & x"e76" => data <= x"0d";
            when "00" & x"e77" => data <= x"11";
            when "00" & x"e78" => data <= x"29";
            when "00" & x"e79" => data <= x"03";
            when "00" & x"e7a" => data <= x"d0";
            when "00" & x"e7b" => data <= x"14";
            when "00" & x"e7c" => data <= x"8a";
            when "00" & x"e7d" => data <= x"d9";
            when "00" & x"e7e" => data <= x"0f";
            when "00" & x"e7f" => data <= x"11";
            when "00" & x"e80" => data <= x"d0";
            when "00" & x"e81" => data <= x"0e";
            when "00" & x"e82" => data <= x"60";
            when "00" & x"e83" => data <= x"b9";
            when "00" & x"e84" => data <= x"0e";
            when "00" & x"e85" => data <= x"11";
            when "00" & x"e86" => data <= x"29";
            when "00" & x"e87" => data <= x"7f";
            when "00" & x"e88" => data <= x"85";
            when "00" & x"e89" => data <= x"ce";
            when "00" & x"e8a" => data <= x"b9";
            when "00" & x"e8b" => data <= x"17";
            when "00" & x"e8c" => data <= x"11";
            when "00" & x"e8d" => data <= x"4c";
            when "00" & x"e8e" => data <= x"7e";
            when "00" & x"e8f" => data <= x"87";
            when "00" & x"e90" => data <= x"4c";
            when "00" & x"e91" => data <= x"af";
            when "00" & x"e92" => data <= x"81";
            when "00" & x"e93" => data <= x"c9";
            when "00" & x"e94" => data <= x"00";
            when "00" & x"e95" => data <= x"d0";
            when "00" & x"e96" => data <= x"06";
            when "00" & x"e97" => data <= x"20";
            when "00" & x"e98" => data <= x"e1";
            when "00" & x"e99" => data <= x"83";
            when "00" & x"e9a" => data <= x"4c";
            when "00" & x"e9b" => data <= x"fa";
            when "00" & x"e9c" => data <= x"8d";
            when "00" & x"e9d" => data <= x"20";
            when "00" & x"e9e" => data <= x"11";
            when "00" & x"e9f" => data <= x"84";
            when "00" & x"ea0" => data <= x"86";
            when "00" & x"ea1" => data <= x"bc";
            when "00" & x"ea2" => data <= x"84";
            when "00" & x"ea3" => data <= x"bd";
            when "00" & x"ea4" => data <= x"85";
            when "00" & x"ea5" => data <= x"b4";
            when "00" & x"ea6" => data <= x"24";
            when "00" & x"ea7" => data <= x"b4";
            when "00" & x"ea8" => data <= x"08";
            when "00" & x"ea9" => data <= x"20";
            when "00" & x"eaa" => data <= x"06";
            when "00" & x"eab" => data <= x"81";
            when "00" & x"eac" => data <= x"20";
            when "00" & x"ead" => data <= x"96";
            when "00" & x"eae" => data <= x"82";
            when "00" & x"eaf" => data <= x"b0";
            when "00" & x"eb0" => data <= x"1a";
            when "00" & x"eb1" => data <= x"28";
            when "00" & x"eb2" => data <= x"50";
            when "00" & x"eb3" => data <= x"03";
            when "00" & x"eb4" => data <= x"a9";
            when "00" & x"eb5" => data <= x"00";
            when "00" & x"eb6" => data <= x"60";
            when "00" & x"eb7" => data <= x"08";
            when "00" & x"eb8" => data <= x"a9";
            when "00" & x"eb9" => data <= x"00";
            when "00" & x"eba" => data <= x"a2";
            when "00" & x"ebb" => data <= x"07";
            when "00" & x"ebc" => data <= x"95";
            when "00" & x"ebd" => data <= x"be";
            when "00" & x"ebe" => data <= x"9d";
            when "00" & x"ebf" => data <= x"74";
            when "00" & x"ec0" => data <= x"10";
            when "00" & x"ec1" => data <= x"ca";
            when "00" & x"ec2" => data <= x"10";
            when "00" & x"ec3" => data <= x"f8";
            when "00" & x"ec4" => data <= x"a9";
            when "00" & x"ec5" => data <= x"40";
            when "00" & x"ec6" => data <= x"85";
            when "00" & x"ec7" => data <= x"c5";
            when "00" & x"ec8" => data <= x"20";
            when "00" & x"ec9" => data <= x"61";
            when "00" & x"eca" => data <= x"89";
            when "00" & x"ecb" => data <= x"28";
            when "00" & x"ecc" => data <= x"08";
            when "00" & x"ecd" => data <= x"70";
            when "00" & x"ece" => data <= x"03";
            when "00" & x"ecf" => data <= x"20";
            when "00" & x"ed0" => data <= x"3c";
            when "00" & x"ed1" => data <= x"98";
            when "00" & x"ed2" => data <= x"20";
            when "00" & x"ed3" => data <= x"9e";
            when "00" & x"ed4" => data <= x"8f";
            when "00" & x"ed5" => data <= x"90";
            when "00" & x"ed6" => data <= x"0e";
            when "00" & x"ed7" => data <= x"b9";
            when "00" & x"ed8" => data <= x"0c";
            when "00" & x"ed9" => data <= x"11";
            when "00" & x"eda" => data <= x"10";
            when "00" & x"edb" => data <= x"26";
            when "00" & x"edc" => data <= x"24";
            when "00" & x"edd" => data <= x"b4";
            when "00" & x"ede" => data <= x"30";
            when "00" & x"edf" => data <= x"22";
            when "00" & x"ee0" => data <= x"20";
            when "00" & x"ee1" => data <= x"99";
            when "00" & x"ee2" => data <= x"8f";
            when "00" & x"ee3" => data <= x"b0";
            when "00" & x"ee4" => data <= x"f2";
            when "00" & x"ee5" => data <= x"ac";
            when "00" & x"ee6" => data <= x"c2";
            when "00" & x"ee7" => data <= x"10";
            when "00" & x"ee8" => data <= x"d0";
            when "00" & x"ee9" => data <= x"21";
            when "00" & x"eea" => data <= x"20";
            when "00" & x"eeb" => data <= x"33";
            when "00" & x"eec" => data <= x"80";
            when "00" & x"eed" => data <= x"c0";
            when "00" & x"eee" => data <= x"54";
            when "00" & x"eef" => data <= x"6f";
            when "00" & x"ef0" => data <= x"6f";
            when "00" & x"ef1" => data <= x"20";
            when "00" & x"ef2" => data <= x"6d";
            when "00" & x"ef3" => data <= x"61";
            when "00" & x"ef4" => data <= x"6e";
            when "00" & x"ef5" => data <= x"79";
            when "00" & x"ef6" => data <= x"20";
            when "00" & x"ef7" => data <= x"66";
            when "00" & x"ef8" => data <= x"69";
            when "00" & x"ef9" => data <= x"6c";
            when "00" & x"efa" => data <= x"65";
            when "00" & x"efb" => data <= x"73";
            when "00" & x"efc" => data <= x"20";
            when "00" & x"efd" => data <= x"6f";
            when "00" & x"efe" => data <= x"70";
            when "00" & x"eff" => data <= x"65";
            when "00" & x"f00" => data <= x"6e";
            when "00" & x"f01" => data <= x"00";
            when "00" & x"f02" => data <= x"20";
            when "00" & x"f03" => data <= x"2b";
            when "00" & x"f04" => data <= x"80";
            when "00" & x"f05" => data <= x"c2";
            when "00" & x"f06" => data <= x"6f";
            when "00" & x"f07" => data <= x"70";
            when "00" & x"f08" => data <= x"65";
            when "00" & x"f09" => data <= x"6e";
            when "00" & x"f0a" => data <= x"00";
            when "00" & x"f0b" => data <= x"a9";
            when "00" & x"f0c" => data <= x"08";
            when "00" & x"f0d" => data <= x"8d";
            when "00" & x"f0e" => data <= x"c5";
            when "00" & x"f0f" => data <= x"10";
            when "00" & x"f10" => data <= x"bd";
            when "00" & x"f11" => data <= x"08";
            when "00" & x"f12" => data <= x"0e";
            when "00" & x"f13" => data <= x"99";
            when "00" & x"f14" => data <= x"00";
            when "00" & x"f15" => data <= x"11";
            when "00" & x"f16" => data <= x"c8";
            when "00" & x"f17" => data <= x"bd";
            when "00" & x"f18" => data <= x"08";
            when "00" & x"f19" => data <= x"0f";
            when "00" & x"f1a" => data <= x"99";
            when "00" & x"f1b" => data <= x"00";
            when "00" & x"f1c" => data <= x"11";
            when "00" & x"f1d" => data <= x"c8";
            when "00" & x"f1e" => data <= x"e8";
            when "00" & x"f1f" => data <= x"ce";
            when "00" & x"f20" => data <= x"c5";
            when "00" & x"f21" => data <= x"10";
            when "00" & x"f22" => data <= x"d0";
            when "00" & x"f23" => data <= x"ec";
            when "00" & x"f24" => data <= x"a2";
            when "00" & x"f25" => data <= x"10";
            when "00" & x"f26" => data <= x"a9";
            when "00" & x"f27" => data <= x"00";
            when "00" & x"f28" => data <= x"99";
            when "00" & x"f29" => data <= x"00";
            when "00" & x"f2a" => data <= x"11";
            when "00" & x"f2b" => data <= x"c8";
            when "00" & x"f2c" => data <= x"ca";
            when "00" & x"f2d" => data <= x"d0";
            when "00" & x"f2e" => data <= x"f9";
            when "00" & x"f2f" => data <= x"ad";
            when "00" & x"f30" => data <= x"c2";
            when "00" & x"f31" => data <= x"10";
            when "00" & x"f32" => data <= x"a8";
            when "00" & x"f33" => data <= x"20";
            when "00" & x"f34" => data <= x"04";
            when "00" & x"f35" => data <= x"82";
            when "00" & x"f36" => data <= x"69";
            when "00" & x"f37" => data <= x"11";
            when "00" & x"f38" => data <= x"99";
            when "00" & x"f39" => data <= x"13";
            when "00" & x"f3a" => data <= x"11";
            when "00" & x"f3b" => data <= x"ad";
            when "00" & x"f3c" => data <= x"c1";
            when "00" & x"f3d" => data <= x"10";
            when "00" & x"f3e" => data <= x"99";
            when "00" & x"f3f" => data <= x"1b";
            when "00" & x"f40" => data <= x"11";
            when "00" & x"f41" => data <= x"0d";
            when "00" & x"f42" => data <= x"c0";
            when "00" & x"f43" => data <= x"10";
            when "00" & x"f44" => data <= x"8d";
            when "00" & x"f45" => data <= x"c0";
            when "00" & x"f46" => data <= x"10";
            when "00" & x"f47" => data <= x"b9";
            when "00" & x"f48" => data <= x"09";
            when "00" & x"f49" => data <= x"11";
            when "00" & x"f4a" => data <= x"69";
            when "00" & x"f4b" => data <= x"ff";
            when "00" & x"f4c" => data <= x"b9";
            when "00" & x"f4d" => data <= x"0b";
            when "00" & x"f4e" => data <= x"11";
            when "00" & x"f4f" => data <= x"69";
            when "00" & x"f50" => data <= x"00";
            when "00" & x"f51" => data <= x"99";
            when "00" & x"f52" => data <= x"19";
            when "00" & x"f53" => data <= x"11";
            when "00" & x"f54" => data <= x"b9";
            when "00" & x"f55" => data <= x"0d";
            when "00" & x"f56" => data <= x"11";
            when "00" & x"f57" => data <= x"09";
            when "00" & x"f58" => data <= x"0f";
            when "00" & x"f59" => data <= x"69";
            when "00" & x"f5a" => data <= x"00";
            when "00" & x"f5b" => data <= x"20";
            when "00" & x"f5c" => data <= x"fd";
            when "00" & x"f5d" => data <= x"81";
            when "00" & x"f5e" => data <= x"99";
            when "00" & x"f5f" => data <= x"1a";
            when "00" & x"f60" => data <= x"11";
            when "00" & x"f61" => data <= x"28";
            when "00" & x"f62" => data <= x"50";
            when "00" & x"f63" => data <= x"2e";
            when "00" & x"f64" => data <= x"30";
            when "00" & x"f65" => data <= x"08";
            when "00" & x"f66" => data <= x"a9";
            when "00" & x"f67" => data <= x"80";
            when "00" & x"f68" => data <= x"19";
            when "00" & x"f69" => data <= x"0c";
            when "00" & x"f6a" => data <= x"11";
            when "00" & x"f6b" => data <= x"99";
            when "00" & x"f6c" => data <= x"0c";
            when "00" & x"f6d" => data <= x"11";
            when "00" & x"f6e" => data <= x"b9";
            when "00" & x"f6f" => data <= x"09";
            when "00" & x"f70" => data <= x"11";
            when "00" & x"f71" => data <= x"99";
            when "00" & x"f72" => data <= x"14";
            when "00" & x"f73" => data <= x"11";
            when "00" & x"f74" => data <= x"b9";
            when "00" & x"f75" => data <= x"0b";
            when "00" & x"f76" => data <= x"11";
            when "00" & x"f77" => data <= x"99";
            when "00" & x"f78" => data <= x"15";
            when "00" & x"f79" => data <= x"11";
            when "00" & x"f7a" => data <= x"b9";
            when "00" & x"f7b" => data <= x"0d";
            when "00" & x"f7c" => data <= x"11";
            when "00" & x"f7d" => data <= x"20";
            when "00" & x"f7e" => data <= x"fd";
            when "00" & x"f7f" => data <= x"81";
            when "00" & x"f80" => data <= x"99";
            when "00" & x"f81" => data <= x"16";
            when "00" & x"f82" => data <= x"11";
            when "00" & x"f83" => data <= x"a5";
            when "00" & x"f84" => data <= x"cf";
            when "00" & x"f85" => data <= x"19";
            when "00" & x"f86" => data <= x"17";
            when "00" & x"f87" => data <= x"11";
            when "00" & x"f88" => data <= x"99";
            when "00" & x"f89" => data <= x"17";
            when "00" & x"f8a" => data <= x"11";
            when "00" & x"f8b" => data <= x"98";
            when "00" & x"f8c" => data <= x"20";
            when "00" & x"f8d" => data <= x"04";
            when "00" & x"f8e" => data <= x"82";
            when "00" & x"f8f" => data <= x"09";
            when "00" & x"f90" => data <= x"10";
            when "00" & x"f91" => data <= x"60";
            when "00" & x"f92" => data <= x"a9";
            when "00" & x"f93" => data <= x"20";
            when "00" & x"f94" => data <= x"99";
            when "00" & x"f95" => data <= x"17";
            when "00" & x"f96" => data <= x"11";
            when "00" & x"f97" => data <= x"d0";
            when "00" & x"f98" => data <= x"ea";
            when "00" & x"f99" => data <= x"8a";
            when "00" & x"f9a" => data <= x"48";
            when "00" & x"f9b" => data <= x"4c";
            when "00" & x"f9c" => data <= x"dd";
            when "00" & x"f9d" => data <= x"8f";
            when "00" & x"f9e" => data <= x"a9";
            when "00" & x"f9f" => data <= x"00";
            when "00" & x"fa0" => data <= x"8d";
            when "00" & x"fa1" => data <= x"c2";
            when "00" & x"fa2" => data <= x"10";
            when "00" & x"fa3" => data <= x"a9";
            when "00" & x"fa4" => data <= x"08";
            when "00" & x"fa5" => data <= x"85";
            when "00" & x"fa6" => data <= x"b5";
            when "00" & x"fa7" => data <= x"98";
            when "00" & x"fa8" => data <= x"aa";
            when "00" & x"fa9" => data <= x"a0";
            when "00" & x"faa" => data <= x"a0";
            when "00" & x"fab" => data <= x"84";
            when "00" & x"fac" => data <= x"b3";
            when "00" & x"fad" => data <= x"8a";
            when "00" & x"fae" => data <= x"48";
            when "00" & x"faf" => data <= x"a9";
            when "00" & x"fb0" => data <= x"08";
            when "00" & x"fb1" => data <= x"85";
            when "00" & x"fb2" => data <= x"b2";
            when "00" & x"fb3" => data <= x"a5";
            when "00" & x"fb4" => data <= x"b5";
            when "00" & x"fb5" => data <= x"2c";
            when "00" & x"fb6" => data <= x"c0";
            when "00" & x"fb7" => data <= x"10";
            when "00" & x"fb8" => data <= x"f0";
            when "00" & x"fb9" => data <= x"1d";
            when "00" & x"fba" => data <= x"b9";
            when "00" & x"fbb" => data <= x"17";
            when "00" & x"fbc" => data <= x"11";
            when "00" & x"fbd" => data <= x"45";
            when "00" & x"fbe" => data <= x"cf";
            when "00" & x"fbf" => data <= x"29";
            when "00" & x"fc0" => data <= x"03";
            when "00" & x"fc1" => data <= x"d0";
            when "00" & x"fc2" => data <= x"1a";
            when "00" & x"fc3" => data <= x"bd";
            when "00" & x"fc4" => data <= x"08";
            when "00" & x"fc5" => data <= x"0e";
            when "00" & x"fc6" => data <= x"59";
            when "00" & x"fc7" => data <= x"00";
            when "00" & x"fc8" => data <= x"11";
            when "00" & x"fc9" => data <= x"29";
            when "00" & x"fca" => data <= x"7f";
            when "00" & x"fcb" => data <= x"d0";
            when "00" & x"fcc" => data <= x"10";
            when "00" & x"fcd" => data <= x"e8";
            when "00" & x"fce" => data <= x"c8";
            when "00" & x"fcf" => data <= x"c8";
            when "00" & x"fd0" => data <= x"c6";
            when "00" & x"fd1" => data <= x"b2";
            when "00" & x"fd2" => data <= x"d0";
            when "00" & x"fd3" => data <= x"ef";
            when "00" & x"fd4" => data <= x"38";
            when "00" & x"fd5" => data <= x"b0";
            when "00" & x"fd6" => data <= x"10";
            when "00" & x"fd7" => data <= x"8c";
            when "00" & x"fd8" => data <= x"c2";
            when "00" & x"fd9" => data <= x"10";
            when "00" & x"fda" => data <= x"8d";
            when "00" & x"fdb" => data <= x"c1";
            when "00" & x"fdc" => data <= x"10";
            when "00" & x"fdd" => data <= x"38";
            when "00" & x"fde" => data <= x"a5";
            when "00" & x"fdf" => data <= x"b3";
            when "00" & x"fe0" => data <= x"e9";
            when "00" & x"fe1" => data <= x"20";
            when "00" & x"fe2" => data <= x"85";
            when "00" & x"fe3" => data <= x"b3";
            when "00" & x"fe4" => data <= x"06";
            when "00" & x"fe5" => data <= x"b5";
            when "00" & x"fe6" => data <= x"18";
            when "00" & x"fe7" => data <= x"68";
            when "00" & x"fe8" => data <= x"aa";
            when "00" & x"fe9" => data <= x"a4";
            when "00" & x"fea" => data <= x"b3";
            when "00" & x"feb" => data <= x"a5";
            when "00" & x"fec" => data <= x"b5";
            when "00" & x"fed" => data <= x"b0";
            when "00" & x"fee" => data <= x"02";
            when "00" & x"fef" => data <= x"d0";
            when "00" & x"ff0" => data <= x"ba";
            when "00" & x"ff1" => data <= x"60";
            when "00" & x"ff2" => data <= x"ad";
            when "00" & x"ff3" => data <= x"c0";
            when "00" & x"ff4" => data <= x"10";
            when "00" & x"ff5" => data <= x"48";
            when "00" & x"ff6" => data <= x"20";
            when "00" & x"ff7" => data <= x"ed";
            when "00" & x"ff8" => data <= x"8d";
            when "00" & x"ff9" => data <= x"f0";
            when "00" & x"ffa" => data <= x"07";
            when "00" & x"ffb" => data <= x"ad";
            when "00" & x"ffc" => data <= x"c0";
            when "00" & x"ffd" => data <= x"10";
            when "00" & x"ffe" => data <= x"48";
            when "00" & x"fff" => data <= x"20";
            when "01" & x"000" => data <= x"fa";
            when "01" & x"001" => data <= x"8d";
            when "01" & x"002" => data <= x"68";
            when "01" & x"003" => data <= x"8d";
            when "01" & x"004" => data <= x"c0";
            when "01" & x"005" => data <= x"10";
            when "01" & x"006" => data <= x"60";
            when "01" & x"007" => data <= x"c0";
            when "01" & x"008" => data <= x"00";
            when "01" & x"009" => data <= x"f0";
            when "01" & x"00a" => data <= x"11";
            when "01" & x"00b" => data <= x"20";
            when "01" & x"00c" => data <= x"e1";
            when "01" & x"00d" => data <= x"83";
            when "01" & x"00e" => data <= x"c9";
            when "01" & x"00f" => data <= x"ff";
            when "01" & x"010" => data <= x"f0";
            when "01" & x"011" => data <= x"e9";
            when "01" & x"012" => data <= x"c9";
            when "01" & x"013" => data <= x"03";
            when "01" & x"014" => data <= x"b0";
            when "01" & x"015" => data <= x"17";
            when "01" & x"016" => data <= x"4a";
            when "01" & x"017" => data <= x"90";
            when "01" & x"018" => data <= x"15";
            when "01" & x"019" => data <= x"4c";
            when "01" & x"01a" => data <= x"a7";
            when "01" & x"01b" => data <= x"92";
            when "01" & x"01c" => data <= x"20";
            when "01" & x"01d" => data <= x"11";
            when "01" & x"01e" => data <= x"84";
            when "01" & x"01f" => data <= x"a8";
            when "01" & x"020" => data <= x"c8";
            when "01" & x"021" => data <= x"c0";
            when "01" & x"022" => data <= x"03";
            when "01" & x"023" => data <= x"b0";
            when "01" & x"024" => data <= x"08";
            when "01" & x"025" => data <= x"b9";
            when "01" & x"026" => data <= x"81";
            when "01" & x"027" => data <= x"99";
            when "01" & x"028" => data <= x"48";
            when "01" & x"029" => data <= x"b9";
            when "01" & x"02a" => data <= x"7e";
            when "01" & x"02b" => data <= x"99";
            when "01" & x"02c" => data <= x"48";
            when "01" & x"02d" => data <= x"60";
            when "01" & x"02e" => data <= x"20";
            when "01" & x"02f" => data <= x"e1";
            when "01" & x"030" => data <= x"83";
            when "01" & x"031" => data <= x"20";
            when "01" & x"032" => data <= x"a5";
            when "01" & x"033" => data <= x"90";
            when "01" & x"034" => data <= x"8c";
            when "01" & x"035" => data <= x"c2";
            when "01" & x"036" => data <= x"10";
            when "01" & x"037" => data <= x"0a";
            when "01" & x"038" => data <= x"0a";
            when "01" & x"039" => data <= x"6d";
            when "01" & x"03a" => data <= x"c2";
            when "01" & x"03b" => data <= x"10";
            when "01" & x"03c" => data <= x"a8";
            when "01" & x"03d" => data <= x"b9";
            when "01" & x"03e" => data <= x"10";
            when "01" & x"03f" => data <= x"11";
            when "01" & x"040" => data <= x"95";
            when "01" & x"041" => data <= x"00";
            when "01" & x"042" => data <= x"b9";
            when "01" & x"043" => data <= x"11";
            when "01" & x"044" => data <= x"11";
            when "01" & x"045" => data <= x"95";
            when "01" & x"046" => data <= x"01";
            when "01" & x"047" => data <= x"b9";
            when "01" & x"048" => data <= x"12";
            when "01" & x"049" => data <= x"11";
            when "01" & x"04a" => data <= x"95";
            when "01" & x"04b" => data <= x"02";
            when "01" & x"04c" => data <= x"a9";
            when "01" & x"04d" => data <= x"00";
            when "01" & x"04e" => data <= x"95";
            when "01" & x"04f" => data <= x"03";
            when "01" & x"050" => data <= x"60";
            when "01" & x"051" => data <= x"48";
            when "01" & x"052" => data <= x"8e";
            when "01" & x"053" => data <= x"c6";
            when "01" & x"054" => data <= x"10";
            when "01" & x"055" => data <= x"98";
            when "01" & x"056" => data <= x"29";
            when "01" & x"057" => data <= x"e0";
            when "01" & x"058" => data <= x"8d";
            when "01" & x"059" => data <= x"c2";
            when "01" & x"05a" => data <= x"10";
            when "01" & x"05b" => data <= x"f0";
            when "01" & x"05c" => data <= x"13";
            when "01" & x"05d" => data <= x"20";
            when "01" & x"05e" => data <= x"04";
            when "01" & x"05f" => data <= x"82";
            when "01" & x"060" => data <= x"a8";
            when "01" & x"061" => data <= x"a9";
            when "01" & x"062" => data <= x"00";
            when "01" & x"063" => data <= x"38";
            when "01" & x"064" => data <= x"6a";
            when "01" & x"065" => data <= x"88";
            when "01" & x"066" => data <= x"d0";
            when "01" & x"067" => data <= x"fc";
            when "01" & x"068" => data <= x"ac";
            when "01" & x"069" => data <= x"c2";
            when "01" & x"06a" => data <= x"10";
            when "01" & x"06b" => data <= x"2c";
            when "01" & x"06c" => data <= x"c0";
            when "01" & x"06d" => data <= x"10";
            when "01" & x"06e" => data <= x"d0";
            when "01" & x"06f" => data <= x"03";
            when "01" & x"070" => data <= x"68";
            when "01" & x"071" => data <= x"38";
            when "01" & x"072" => data <= x"60";
            when "01" & x"073" => data <= x"68";
            when "01" & x"074" => data <= x"18";
            when "01" & x"075" => data <= x"60";
            when "01" & x"076" => data <= x"48";
            when "01" & x"077" => data <= x"8a";
            when "01" & x"078" => data <= x"4c";
            when "01" & x"079" => data <= x"7d";
            when "01" & x"07a" => data <= x"90";
            when "01" & x"07b" => data <= x"48";
            when "01" & x"07c" => data <= x"98";
            when "01" & x"07d" => data <= x"c9";
            when "01" & x"07e" => data <= x"10";
            when "01" & x"07f" => data <= x"90";
            when "01" & x"080" => data <= x"04";
            when "01" & x"081" => data <= x"c9";
            when "01" & x"082" => data <= x"18";
            when "01" & x"083" => data <= x"90";
            when "01" & x"084" => data <= x"02";
            when "01" & x"085" => data <= x"a9";
            when "01" & x"086" => data <= x"08";
            when "01" & x"087" => data <= x"20";
            when "01" & x"088" => data <= x"0a";
            when "01" & x"089" => data <= x"82";
            when "01" & x"08a" => data <= x"a8";
            when "01" & x"08b" => data <= x"68";
            when "01" & x"08c" => data <= x"60";
            when "01" & x"08d" => data <= x"48";
            when "01" & x"08e" => data <= x"98";
            when "01" & x"08f" => data <= x"48";
            when "01" & x"090" => data <= x"8a";
            when "01" & x"091" => data <= x"a8";
            when "01" & x"092" => data <= x"20";
            when "01" & x"093" => data <= x"a5";
            when "01" & x"094" => data <= x"90";
            when "01" & x"095" => data <= x"98";
            when "01" & x"096" => data <= x"20";
            when "01" & x"097" => data <= x"f8";
            when "01" & x"098" => data <= x"92";
            when "01" & x"099" => data <= x"d0";
            when "01" & x"09a" => data <= x"04";
            when "01" & x"09b" => data <= x"a2";
            when "01" & x"09c" => data <= x"ff";
            when "01" & x"09d" => data <= x"d0";
            when "01" & x"09e" => data <= x"02";
            when "01" & x"09f" => data <= x"a2";
            when "01" & x"0a0" => data <= x"00";
            when "01" & x"0a1" => data <= x"68";
            when "01" & x"0a2" => data <= x"a8";
            when "01" & x"0a3" => data <= x"68";
            when "01" & x"0a4" => data <= x"60";
            when "01" & x"0a5" => data <= x"20";
            when "01" & x"0a6" => data <= x"7b";
            when "01" & x"0a7" => data <= x"90";
            when "01" & x"0a8" => data <= x"20";
            when "01" & x"0a9" => data <= x"51";
            when "01" & x"0aa" => data <= x"90";
            when "01" & x"0ab" => data <= x"90";
            when "01" & x"0ac" => data <= x"f7";
            when "01" & x"0ad" => data <= x"20";
            when "01" & x"0ae" => data <= x"33";
            when "01" & x"0af" => data <= x"80";
            when "01" & x"0b0" => data <= x"de";
            when "01" & x"0b1" => data <= x"43";
            when "01" & x"0b2" => data <= x"68";
            when "01" & x"0b3" => data <= x"61";
            when "01" & x"0b4" => data <= x"6e";
            when "01" & x"0b5" => data <= x"6e";
            when "01" & x"0b6" => data <= x"65";
            when "01" & x"0b7" => data <= x"6c";
            when "01" & x"0b8" => data <= x"00";
            when "01" & x"0b9" => data <= x"20";
            when "01" & x"0ba" => data <= x"33";
            when "01" & x"0bb" => data <= x"80";
            when "01" & x"0bc" => data <= x"df";
            when "01" & x"0bd" => data <= x"45";
            when "01" & x"0be" => data <= x"4f";
            when "01" & x"0bf" => data <= x"46";
            when "01" & x"0c0" => data <= x"00";
            when "01" & x"0c1" => data <= x"20";
            when "01" & x"0c2" => data <= x"11";
            when "01" & x"0c3" => data <= x"84";
            when "01" & x"0c4" => data <= x"20";
            when "01" & x"0c5" => data <= x"a5";
            when "01" & x"0c6" => data <= x"90";
            when "01" & x"0c7" => data <= x"98";
            when "01" & x"0c8" => data <= x"20";
            when "01" & x"0c9" => data <= x"f8";
            when "01" & x"0ca" => data <= x"92";
            when "01" & x"0cb" => data <= x"d0";
            when "01" & x"0cc" => data <= x"13";
            when "01" & x"0cd" => data <= x"b9";
            when "01" & x"0ce" => data <= x"17";
            when "01" & x"0cf" => data <= x"11";
            when "01" & x"0d0" => data <= x"29";
            when "01" & x"0d1" => data <= x"10";
            when "01" & x"0d2" => data <= x"d0";
            when "01" & x"0d3" => data <= x"e5";
            when "01" & x"0d4" => data <= x"a9";
            when "01" & x"0d5" => data <= x"10";
            when "01" & x"0d6" => data <= x"20";
            when "01" & x"0d7" => data <= x"3c";
            when "01" & x"0d8" => data <= x"91";
            when "01" & x"0d9" => data <= x"ae";
            when "01" & x"0da" => data <= x"c6";
            when "01" & x"0db" => data <= x"10";
            when "01" & x"0dc" => data <= x"a9";
            when "01" & x"0dd" => data <= x"fe";
            when "01" & x"0de" => data <= x"38";
            when "01" & x"0df" => data <= x"60";
            when "01" & x"0e0" => data <= x"b9";
            when "01" & x"0e1" => data <= x"17";
            when "01" & x"0e2" => data <= x"11";
            when "01" & x"0e3" => data <= x"30";
            when "01" & x"0e4" => data <= x"0a";
            when "01" & x"0e5" => data <= x"20";
            when "01" & x"0e6" => data <= x"83";
            when "01" & x"0e7" => data <= x"8e";
            when "01" & x"0e8" => data <= x"20";
            when "01" & x"0e9" => data <= x"4b";
            when "01" & x"0ea" => data <= x"91";
            when "01" & x"0eb" => data <= x"38";
            when "01" & x"0ec" => data <= x"20";
            when "01" & x"0ed" => data <= x"53";
            when "01" & x"0ee" => data <= x"91";
            when "01" & x"0ef" => data <= x"b9";
            when "01" & x"0f0" => data <= x"10";
            when "01" & x"0f1" => data <= x"11";
            when "01" & x"0f2" => data <= x"85";
            when "01" & x"0f3" => data <= x"bc";
            when "01" & x"0f4" => data <= x"b9";
            when "01" & x"0f5" => data <= x"13";
            when "01" & x"0f6" => data <= x"11";
            when "01" & x"0f7" => data <= x"85";
            when "01" & x"0f8" => data <= x"bd";
            when "01" & x"0f9" => data <= x"a0";
            when "01" & x"0fa" => data <= x"00";
            when "01" & x"0fb" => data <= x"b1";
            when "01" & x"0fc" => data <= x"bc";
            when "01" & x"0fd" => data <= x"48";
            when "01" & x"0fe" => data <= x"ac";
            when "01" & x"0ff" => data <= x"c2";
            when "01" & x"100" => data <= x"10";
            when "01" & x"101" => data <= x"a6";
            when "01" & x"102" => data <= x"bc";
            when "01" & x"103" => data <= x"e8";
            when "01" & x"104" => data <= x"8a";
            when "01" & x"105" => data <= x"99";
            when "01" & x"106" => data <= x"10";
            when "01" & x"107" => data <= x"11";
            when "01" & x"108" => data <= x"d0";
            when "01" & x"109" => data <= x"14";
            when "01" & x"10a" => data <= x"18";
            when "01" & x"10b" => data <= x"b9";
            when "01" & x"10c" => data <= x"11";
            when "01" & x"10d" => data <= x"11";
            when "01" & x"10e" => data <= x"69";
            when "01" & x"10f" => data <= x"01";
            when "01" & x"110" => data <= x"99";
            when "01" & x"111" => data <= x"11";
            when "01" & x"112" => data <= x"11";
            when "01" & x"113" => data <= x"b9";
            when "01" & x"114" => data <= x"12";
            when "01" & x"115" => data <= x"11";
            when "01" & x"116" => data <= x"69";
            when "01" & x"117" => data <= x"00";
            when "01" & x"118" => data <= x"99";
            when "01" & x"119" => data <= x"12";
            when "01" & x"11a" => data <= x"11";
            when "01" & x"11b" => data <= x"20";
            when "01" & x"11c" => data <= x"41";
            when "01" & x"11d" => data <= x"91";
            when "01" & x"11e" => data <= x"18";
            when "01" & x"11f" => data <= x"68";
            when "01" & x"120" => data <= x"60";
            when "01" & x"121" => data <= x"18";
            when "01" & x"122" => data <= x"b9";
            when "01" & x"123" => data <= x"0f";
            when "01" & x"124" => data <= x"11";
            when "01" & x"125" => data <= x"79";
            when "01" & x"126" => data <= x"11";
            when "01" & x"127" => data <= x"11";
            when "01" & x"128" => data <= x"85";
            when "01" & x"129" => data <= x"c5";
            when "01" & x"12a" => data <= x"99";
            when "01" & x"12b" => data <= x"1c";
            when "01" & x"12c" => data <= x"11";
            when "01" & x"12d" => data <= x"b9";
            when "01" & x"12e" => data <= x"0d";
            when "01" & x"12f" => data <= x"11";
            when "01" & x"130" => data <= x"29";
            when "01" & x"131" => data <= x"03";
            when "01" & x"132" => data <= x"79";
            when "01" & x"133" => data <= x"12";
            when "01" & x"134" => data <= x"11";
            when "01" & x"135" => data <= x"85";
            when "01" & x"136" => data <= x"c4";
            when "01" & x"137" => data <= x"99";
            when "01" & x"138" => data <= x"1d";
            when "01" & x"139" => data <= x"11";
            when "01" & x"13a" => data <= x"a9";
            when "01" & x"13b" => data <= x"80";
            when "01" & x"13c" => data <= x"19";
            when "01" & x"13d" => data <= x"17";
            when "01" & x"13e" => data <= x"11";
            when "01" & x"13f" => data <= x"d0";
            when "01" & x"140" => data <= x"05";
            when "01" & x"141" => data <= x"a9";
            when "01" & x"142" => data <= x"7f";
            when "01" & x"143" => data <= x"39";
            when "01" & x"144" => data <= x"17";
            when "01" & x"145" => data <= x"11";
            when "01" & x"146" => data <= x"99";
            when "01" & x"147" => data <= x"17";
            when "01" & x"148" => data <= x"11";
            when "01" & x"149" => data <= x"18";
            when "01" & x"14a" => data <= x"60";
            when "01" & x"14b" => data <= x"b9";
            when "01" & x"14c" => data <= x"17";
            when "01" & x"14d" => data <= x"11";
            when "01" & x"14e" => data <= x"29";
            when "01" & x"14f" => data <= x"40";
            when "01" & x"150" => data <= x"f0";
            when "01" & x"151" => data <= x"3d";
            when "01" & x"152" => data <= x"18";
            when "01" & x"153" => data <= x"08";
            when "01" & x"154" => data <= x"20";
            when "01" & x"155" => data <= x"3e";
            when "01" & x"156" => data <= x"be";
            when "01" & x"157" => data <= x"ac";
            when "01" & x"158" => data <= x"c2";
            when "01" & x"159" => data <= x"10";
            when "01" & x"15a" => data <= x"b9";
            when "01" & x"15b" => data <= x"13";
            when "01" & x"15c" => data <= x"11";
            when "01" & x"15d" => data <= x"85";
            when "01" & x"15e" => data <= x"bf";
            when "01" & x"15f" => data <= x"20";
            when "01" & x"160" => data <= x"8d";
            when "01" & x"161" => data <= x"a0";
            when "01" & x"162" => data <= x"a9";
            when "01" & x"163" => data <= x"00";
            when "01" & x"164" => data <= x"85";
            when "01" & x"165" => data <= x"be";
            when "01" & x"166" => data <= x"85";
            when "01" & x"167" => data <= x"c2";
            when "01" & x"168" => data <= x"a9";
            when "01" & x"169" => data <= x"01";
            when "01" & x"16a" => data <= x"85";
            when "01" & x"16b" => data <= x"c3";
            when "01" & x"16c" => data <= x"28";
            when "01" & x"16d" => data <= x"b0";
            when "01" & x"16e" => data <= x"17";
            when "01" & x"16f" => data <= x"b9";
            when "01" & x"170" => data <= x"1c";
            when "01" & x"171" => data <= x"11";
            when "01" & x"172" => data <= x"85";
            when "01" & x"173" => data <= x"c5";
            when "01" & x"174" => data <= x"b9";
            when "01" & x"175" => data <= x"1d";
            when "01" & x"176" => data <= x"11";
            when "01" & x"177" => data <= x"85";
            when "01" & x"178" => data <= x"c4";
            when "01" & x"179" => data <= x"20";
            when "01" & x"17a" => data <= x"8f";
            when "01" & x"17b" => data <= x"87";
            when "01" & x"17c" => data <= x"ac";
            when "01" & x"17d" => data <= x"c2";
            when "01" & x"17e" => data <= x"10";
            when "01" & x"17f" => data <= x"a9";
            when "01" & x"180" => data <= x"bf";
            when "01" & x"181" => data <= x"20";
            when "01" & x"182" => data <= x"43";
            when "01" & x"183" => data <= x"91";
            when "01" & x"184" => data <= x"90";
            when "01" & x"185" => data <= x"06";
            when "01" & x"186" => data <= x"20";
            when "01" & x"187" => data <= x"21";
            when "01" & x"188" => data <= x"91";
            when "01" & x"189" => data <= x"20";
            when "01" & x"18a" => data <= x"c6";
            when "01" & x"18b" => data <= x"87";
            when "01" & x"18c" => data <= x"ac";
            when "01" & x"18d" => data <= x"c2";
            when "01" & x"18e" => data <= x"10";
            when "01" & x"18f" => data <= x"60";
            when "01" & x"190" => data <= x"4c";
            when "01" & x"191" => data <= x"ad";
            when "01" & x"192" => data <= x"90";
            when "01" & x"193" => data <= x"4c";
            when "01" & x"194" => data <= x"41";
            when "01" & x"195" => data <= x"98";
            when "01" & x"196" => data <= x"20";
            when "01" & x"197" => data <= x"2b";
            when "01" & x"198" => data <= x"80";
            when "01" & x"199" => data <= x"c1";
            when "01" & x"19a" => data <= x"72";
            when "01" & x"19b" => data <= x"65";
            when "01" & x"19c" => data <= x"61";
            when "01" & x"19d" => data <= x"64";
            when "01" & x"19e" => data <= x"20";
            when "01" & x"19f" => data <= x"6f";
            when "01" & x"1a0" => data <= x"6e";
            when "01" & x"1a1" => data <= x"6c";
            when "01" & x"1a2" => data <= x"79";
            when "01" & x"1a3" => data <= x"00";
            when "01" & x"1a4" => data <= x"20";
            when "01" & x"1a5" => data <= x"e1";
            when "01" & x"1a6" => data <= x"83";
            when "01" & x"1a7" => data <= x"4c";
            when "01" & x"1a8" => data <= x"b0";
            when "01" & x"1a9" => data <= x"91";
            when "01" & x"1aa" => data <= x"20";
            when "01" & x"1ab" => data <= x"e1";
            when "01" & x"1ac" => data <= x"83";
            when "01" & x"1ad" => data <= x"20";
            when "01" & x"1ae" => data <= x"a5";
            when "01" & x"1af" => data <= x"90";
            when "01" & x"1b0" => data <= x"48";
            when "01" & x"1b1" => data <= x"b9";
            when "01" & x"1b2" => data <= x"0c";
            when "01" & x"1b3" => data <= x"11";
            when "01" & x"1b4" => data <= x"30";
            when "01" & x"1b5" => data <= x"e0";
            when "01" & x"1b6" => data <= x"b9";
            when "01" & x"1b7" => data <= x"0e";
            when "01" & x"1b8" => data <= x"11";
            when "01" & x"1b9" => data <= x"30";
            when "01" & x"1ba" => data <= x"d8";
            when "01" & x"1bb" => data <= x"20";
            when "01" & x"1bc" => data <= x"83";
            when "01" & x"1bd" => data <= x"8e";
            when "01" & x"1be" => data <= x"98";
            when "01" & x"1bf" => data <= x"18";
            when "01" & x"1c0" => data <= x"69";
            when "01" & x"1c1" => data <= x"04";
            when "01" & x"1c2" => data <= x"20";
            when "01" & x"1c3" => data <= x"f8";
            when "01" & x"1c4" => data <= x"92";
            when "01" & x"1c5" => data <= x"d0";
            when "01" & x"1c6" => data <= x"76";
            when "01" & x"1c7" => data <= x"20";
            when "01" & x"1c8" => data <= x"58";
            when "01" & x"1c9" => data <= x"8e";
            when "01" & x"1ca" => data <= x"ae";
            when "01" & x"1cb" => data <= x"c4";
            when "01" & x"1cc" => data <= x"10";
            when "01" & x"1cd" => data <= x"38";
            when "01" & x"1ce" => data <= x"bd";
            when "01" & x"1cf" => data <= x"07";
            when "01" & x"1d0" => data <= x"0f";
            when "01" & x"1d1" => data <= x"fd";
            when "01" & x"1d2" => data <= x"0f";
            when "01" & x"1d3" => data <= x"0f";
            when "01" & x"1d4" => data <= x"48";
            when "01" & x"1d5" => data <= x"bd";
            when "01" & x"1d6" => data <= x"06";
            when "01" & x"1d7" => data <= x"0f";
            when "01" & x"1d8" => data <= x"fd";
            when "01" & x"1d9" => data <= x"0e";
            when "01" & x"1da" => data <= x"0f";
            when "01" & x"1db" => data <= x"29";
            when "01" & x"1dc" => data <= x"03";
            when "01" & x"1dd" => data <= x"8d";
            when "01" & x"1de" => data <= x"c3";
            when "01" & x"1df" => data <= x"10";
            when "01" & x"1e0" => data <= x"0a";
            when "01" & x"1e1" => data <= x"0a";
            when "01" & x"1e2" => data <= x"0a";
            when "01" & x"1e3" => data <= x"0a";
            when "01" & x"1e4" => data <= x"5d";
            when "01" & x"1e5" => data <= x"0e";
            when "01" & x"1e6" => data <= x"0f";
            when "01" & x"1e7" => data <= x"29";
            when "01" & x"1e8" => data <= x"30";
            when "01" & x"1e9" => data <= x"5d";
            when "01" & x"1ea" => data <= x"0e";
            when "01" & x"1eb" => data <= x"0f";
            when "01" & x"1ec" => data <= x"9d";
            when "01" & x"1ed" => data <= x"0e";
            when "01" & x"1ee" => data <= x"0f";
            when "01" & x"1ef" => data <= x"ad";
            when "01" & x"1f0" => data <= x"c3";
            when "01" & x"1f1" => data <= x"10";
            when "01" & x"1f2" => data <= x"d9";
            when "01" & x"1f3" => data <= x"1a";
            when "01" & x"1f4" => data <= x"11";
            when "01" & x"1f5" => data <= x"d0";
            when "01" & x"1f6" => data <= x"2b";
            when "01" & x"1f7" => data <= x"68";
            when "01" & x"1f8" => data <= x"d9";
            when "01" & x"1f9" => data <= x"19";
            when "01" & x"1fa" => data <= x"11";
            when "01" & x"1fb" => data <= x"d0";
            when "01" & x"1fc" => data <= x"26";
            when "01" & x"1fd" => data <= x"84";
            when "01" & x"1fe" => data <= x"b4";
            when "01" & x"1ff" => data <= x"20";
            when "01" & x"200" => data <= x"20";
            when "01" & x"201" => data <= x"99";
            when "01" & x"202" => data <= x"20";
            when "01" & x"203" => data <= x"76";
            when "01" & x"204" => data <= x"90";
            when "01" & x"205" => data <= x"c4";
            when "01" & x"206" => data <= x"b4";
            when "01" & x"207" => data <= x"d0";
            when "01" & x"208" => data <= x"03";
            when "01" & x"209" => data <= x"20";
            when "01" & x"20a" => data <= x"11";
            when "01" & x"20b" => data <= x"99";
            when "01" & x"20c" => data <= x"a4";
            when "01" & x"20d" => data <= x"b4";
            when "01" & x"20e" => data <= x"20";
            when "01" & x"20f" => data <= x"05";
            when "01" & x"210" => data <= x"8e";
            when "01" & x"211" => data <= x"20";
            when "01" & x"212" => data <= x"33";
            when "01" & x"213" => data <= x"80";
            when "01" & x"214" => data <= x"bf";
            when "01" & x"215" => data <= x"43";
            when "01" & x"216" => data <= x"61";
            when "01" & x"217" => data <= x"6e";
            when "01" & x"218" => data <= x"27";
            when "01" & x"219" => data <= x"74";
            when "01" & x"21a" => data <= x"20";
            when "01" & x"21b" => data <= x"65";
            when "01" & x"21c" => data <= x"78";
            when "01" & x"21d" => data <= x"74";
            when "01" & x"21e" => data <= x"65";
            when "01" & x"21f" => data <= x"6e";
            when "01" & x"220" => data <= x"64";
            when "01" & x"221" => data <= x"00";
            when "01" & x"222" => data <= x"68";
            when "01" & x"223" => data <= x"9d";
            when "01" & x"224" => data <= x"0d";
            when "01" & x"225" => data <= x"0f";
            when "01" & x"226" => data <= x"99";
            when "01" & x"227" => data <= x"19";
            when "01" & x"228" => data <= x"11";
            when "01" & x"229" => data <= x"ad";
            when "01" & x"22a" => data <= x"c3";
            when "01" & x"22b" => data <= x"10";
            when "01" & x"22c" => data <= x"99";
            when "01" & x"22d" => data <= x"1a";
            when "01" & x"22e" => data <= x"11";
            when "01" & x"22f" => data <= x"a9";
            when "01" & x"230" => data <= x"00";
            when "01" & x"231" => data <= x"9d";
            when "01" & x"232" => data <= x"0c";
            when "01" & x"233" => data <= x"0f";
            when "01" & x"234" => data <= x"20";
            when "01" & x"235" => data <= x"b4";
            when "01" & x"236" => data <= x"8a";
            when "01" & x"237" => data <= x"ea";
            when "01" & x"238" => data <= x"ea";
            when "01" & x"239" => data <= x"ea";
            when "01" & x"23a" => data <= x"ac";
            when "01" & x"23b" => data <= x"c2";
            when "01" & x"23c" => data <= x"10";
            when "01" & x"23d" => data <= x"b9";
            when "01" & x"23e" => data <= x"17";
            when "01" & x"23f" => data <= x"11";
            when "01" & x"240" => data <= x"30";
            when "01" & x"241" => data <= x"17";
            when "01" & x"242" => data <= x"20";
            when "01" & x"243" => data <= x"4b";
            when "01" & x"244" => data <= x"91";
            when "01" & x"245" => data <= x"b9";
            when "01" & x"246" => data <= x"14";
            when "01" & x"247" => data <= x"11";
            when "01" & x"248" => data <= x"d0";
            when "01" & x"249" => data <= x"0b";
            when "01" & x"24a" => data <= x"98";
            when "01" & x"24b" => data <= x"20";
            when "01" & x"24c" => data <= x"f8";
            when "01" & x"24d" => data <= x"92";
            when "01" & x"24e" => data <= x"d0";
            when "01" & x"24f" => data <= x"05";
            when "01" & x"250" => data <= x"20";
            when "01" & x"251" => data <= x"21";
            when "01" & x"252" => data <= x"91";
            when "01" & x"253" => data <= x"d0";
            when "01" & x"254" => data <= x"04";
            when "01" & x"255" => data <= x"38";
            when "01" & x"256" => data <= x"20";
            when "01" & x"257" => data <= x"53";
            when "01" & x"258" => data <= x"91";
            when "01" & x"259" => data <= x"b9";
            when "01" & x"25a" => data <= x"10";
            when "01" & x"25b" => data <= x"11";
            when "01" & x"25c" => data <= x"85";
            when "01" & x"25d" => data <= x"bc";
            when "01" & x"25e" => data <= x"b9";
            when "01" & x"25f" => data <= x"13";
            when "01" & x"260" => data <= x"11";
            when "01" & x"261" => data <= x"85";
            when "01" & x"262" => data <= x"bd";
            when "01" & x"263" => data <= x"68";
            when "01" & x"264" => data <= x"a0";
            when "01" & x"265" => data <= x"00";
            when "01" & x"266" => data <= x"91";
            when "01" & x"267" => data <= x"bc";
            when "01" & x"268" => data <= x"ac";
            when "01" & x"269" => data <= x"c2";
            when "01" & x"26a" => data <= x"10";
            when "01" & x"26b" => data <= x"a9";
            when "01" & x"26c" => data <= x"40";
            when "01" & x"26d" => data <= x"20";
            when "01" & x"26e" => data <= x"3c";
            when "01" & x"26f" => data <= x"91";
            when "01" & x"270" => data <= x"e6";
            when "01" & x"271" => data <= x"bc";
            when "01" & x"272" => data <= x"a5";
            when "01" & x"273" => data <= x"bc";
            when "01" & x"274" => data <= x"99";
            when "01" & x"275" => data <= x"10";
            when "01" & x"276" => data <= x"11";
            when "01" & x"277" => data <= x"d0";
            when "01" & x"278" => data <= x"13";
            when "01" & x"279" => data <= x"20";
            when "01" & x"27a" => data <= x"41";
            when "01" & x"27b" => data <= x"91";
            when "01" & x"27c" => data <= x"b9";
            when "01" & x"27d" => data <= x"11";
            when "01" & x"27e" => data <= x"11";
            when "01" & x"27f" => data <= x"69";
            when "01" & x"280" => data <= x"01";
            when "01" & x"281" => data <= x"99";
            when "01" & x"282" => data <= x"11";
            when "01" & x"283" => data <= x"11";
            when "01" & x"284" => data <= x"b9";
            when "01" & x"285" => data <= x"12";
            when "01" & x"286" => data <= x"11";
            when "01" & x"287" => data <= x"69";
            when "01" & x"288" => data <= x"00";
            when "01" & x"289" => data <= x"99";
            when "01" & x"28a" => data <= x"12";
            when "01" & x"28b" => data <= x"11";
            when "01" & x"28c" => data <= x"98";
            when "01" & x"28d" => data <= x"20";
            when "01" & x"28e" => data <= x"f8";
            when "01" & x"28f" => data <= x"92";
            when "01" & x"290" => data <= x"90";
            when "01" & x"291" => data <= x"14";
            when "01" & x"292" => data <= x"a9";
            when "01" & x"293" => data <= x"20";
            when "01" & x"294" => data <= x"20";
            when "01" & x"295" => data <= x"3c";
            when "01" & x"296" => data <= x"91";
            when "01" & x"297" => data <= x"a2";
            when "01" & x"298" => data <= x"02";
            when "01" & x"299" => data <= x"b9";
            when "01" & x"29a" => data <= x"10";
            when "01" & x"29b" => data <= x"11";
            when "01" & x"29c" => data <= x"99";
            when "01" & x"29d" => data <= x"14";
            when "01" & x"29e" => data <= x"11";
            when "01" & x"29f" => data <= x"c8";
            when "01" & x"2a0" => data <= x"ca";
            when "01" & x"2a1" => data <= x"10";
            when "01" & x"2a2" => data <= x"f6";
            when "01" & x"2a3" => data <= x"88";
            when "01" & x"2a4" => data <= x"88";
            when "01" & x"2a5" => data <= x"88";
            when "01" & x"2a6" => data <= x"60";
            when "01" & x"2a7" => data <= x"20";
            when "01" & x"2a8" => data <= x"e1";
            when "01" & x"2a9" => data <= x"83";
            when "01" & x"2aa" => data <= x"20";
            when "01" & x"2ab" => data <= x"a5";
            when "01" & x"2ac" => data <= x"90";
            when "01" & x"2ad" => data <= x"20";
            when "01" & x"2ae" => data <= x"63";
            when "01" & x"2af" => data <= x"a1";
            when "01" & x"2b0" => data <= x"ea";
            when "01" & x"2b1" => data <= x"ea";
            when "01" & x"2b2" => data <= x"ea";
            when "01" & x"2b3" => data <= x"ea";
            when "01" & x"2b4" => data <= x"ea";
            when "01" & x"2b5" => data <= x"ea";
            when "01" & x"2b6" => data <= x"20";
            when "01" & x"2b7" => data <= x"10";
            when "01" & x"2b8" => data <= x"93";
            when "01" & x"2b9" => data <= x"b0";
            when "01" & x"2ba" => data <= x"08";
            when "01" & x"2bb" => data <= x"a9";
            when "01" & x"2bc" => data <= x"00";
            when "01" & x"2bd" => data <= x"20";
            when "01" & x"2be" => data <= x"a4";
            when "01" & x"2bf" => data <= x"91";
            when "01" & x"2c0" => data <= x"4c";
            when "01" & x"2c1" => data <= x"b6";
            when "01" & x"2c2" => data <= x"92";
            when "01" & x"2c3" => data <= x"b5";
            when "01" & x"2c4" => data <= x"00";
            when "01" & x"2c5" => data <= x"99";
            when "01" & x"2c6" => data <= x"10";
            when "01" & x"2c7" => data <= x"11";
            when "01" & x"2c8" => data <= x"b5";
            when "01" & x"2c9" => data <= x"01";
            when "01" & x"2ca" => data <= x"99";
            when "01" & x"2cb" => data <= x"11";
            when "01" & x"2cc" => data <= x"11";
            when "01" & x"2cd" => data <= x"b5";
            when "01" & x"2ce" => data <= x"02";
            when "01" & x"2cf" => data <= x"99";
            when "01" & x"2d0" => data <= x"12";
            when "01" & x"2d1" => data <= x"11";
            when "01" & x"2d2" => data <= x"a9";
            when "01" & x"2d3" => data <= x"6f";
            when "01" & x"2d4" => data <= x"20";
            when "01" & x"2d5" => data <= x"43";
            when "01" & x"2d6" => data <= x"91";
            when "01" & x"2d7" => data <= x"b9";
            when "01" & x"2d8" => data <= x"0f";
            when "01" & x"2d9" => data <= x"11";
            when "01" & x"2da" => data <= x"79";
            when "01" & x"2db" => data <= x"11";
            when "01" & x"2dc" => data <= x"11";
            when "01" & x"2dd" => data <= x"8d";
            when "01" & x"2de" => data <= x"c5";
            when "01" & x"2df" => data <= x"10";
            when "01" & x"2e0" => data <= x"b9";
            when "01" & x"2e1" => data <= x"0d";
            when "01" & x"2e2" => data <= x"11";
            when "01" & x"2e3" => data <= x"29";
            when "01" & x"2e4" => data <= x"03";
            when "01" & x"2e5" => data <= x"79";
            when "01" & x"2e6" => data <= x"12";
            when "01" & x"2e7" => data <= x"11";
            when "01" & x"2e8" => data <= x"d9";
            when "01" & x"2e9" => data <= x"1d";
            when "01" & x"2ea" => data <= x"11";
            when "01" & x"2eb" => data <= x"d0";
            when "01" & x"2ec" => data <= x"b9";
            when "01" & x"2ed" => data <= x"ad";
            when "01" & x"2ee" => data <= x"c5";
            when "01" & x"2ef" => data <= x"10";
            when "01" & x"2f0" => data <= x"d9";
            when "01" & x"2f1" => data <= x"1c";
            when "01" & x"2f2" => data <= x"11";
            when "01" & x"2f3" => data <= x"d0";
            when "01" & x"2f4" => data <= x"b1";
            when "01" & x"2f5" => data <= x"4c";
            when "01" & x"2f6" => data <= x"3a";
            when "01" & x"2f7" => data <= x"91";
            when "01" & x"2f8" => data <= x"aa";
            when "01" & x"2f9" => data <= x"b9";
            when "01" & x"2fa" => data <= x"12";
            when "01" & x"2fb" => data <= x"11";
            when "01" & x"2fc" => data <= x"dd";
            when "01" & x"2fd" => data <= x"16";
            when "01" & x"2fe" => data <= x"11";
            when "01" & x"2ff" => data <= x"d0";
            when "01" & x"300" => data <= x"0e";
            when "01" & x"301" => data <= x"b9";
            when "01" & x"302" => data <= x"11";
            when "01" & x"303" => data <= x"11";
            when "01" & x"304" => data <= x"dd";
            when "01" & x"305" => data <= x"15";
            when "01" & x"306" => data <= x"11";
            when "01" & x"307" => data <= x"d0";
            when "01" & x"308" => data <= x"06";
            when "01" & x"309" => data <= x"b9";
            when "01" & x"30a" => data <= x"10";
            when "01" & x"30b" => data <= x"11";
            when "01" & x"30c" => data <= x"dd";
            when "01" & x"30d" => data <= x"14";
            when "01" & x"30e" => data <= x"11";
            when "01" & x"30f" => data <= x"60";
            when "01" & x"310" => data <= x"b9";
            when "01" & x"311" => data <= x"14";
            when "01" & x"312" => data <= x"11";
            when "01" & x"313" => data <= x"d5";
            when "01" & x"314" => data <= x"00";
            when "01" & x"315" => data <= x"b9";
            when "01" & x"316" => data <= x"15";
            when "01" & x"317" => data <= x"11";
            when "01" & x"318" => data <= x"f5";
            when "01" & x"319" => data <= x"01";
            when "01" & x"31a" => data <= x"b9";
            when "01" & x"31b" => data <= x"16";
            when "01" & x"31c" => data <= x"11";
            when "01" & x"31d" => data <= x"f5";
            when "01" & x"31e" => data <= x"02";
            when "01" & x"31f" => data <= x"60";
            when "01" & x"320" => data <= x"a5";
            when "01" & x"321" => data <= x"b3";
            when "01" & x"322" => data <= x"48";
            when "01" & x"323" => data <= x"a9";
            when "01" & x"324" => data <= x"ff";
            when "01" & x"325" => data <= x"8d";
            when "01" & x"326" => data <= x"de";
            when "01" & x"327" => data <= x"10";
            when "01" & x"328" => data <= x"20";
            when "01" & x"329" => data <= x"65";
            when "01" & x"32a" => data <= x"80";
            when "01" & x"32b" => data <= x"53";
            when "01" & x"32c" => data <= x"6d";
            when "01" & x"32d" => data <= x"61";
            when "01" & x"32e" => data <= x"72";
            when "01" & x"32f" => data <= x"74";
            when "01" & x"330" => data <= x"20";
            when "01" & x"331" => data <= x"53";
            when "01" & x"332" => data <= x"50";
            when "01" & x"333" => data <= x"49";
            when "01" & x"334" => data <= x"0d";
            when "01" & x"335" => data <= x"0d";
            when "01" & x"336" => data <= x"90";
            when "01" & x"337" => data <= x"03";
            when "01" & x"338" => data <= x"4c";
            when "01" & x"339" => data <= x"28";
            when "01" & x"33a" => data <= x"b1";
            when "01" & x"33b" => data <= x"a9";
            when "01" & x"33c" => data <= x"00";
            when "01" & x"33d" => data <= x"ba";
            when "01" & x"33e" => data <= x"9d";
            when "01" & x"33f" => data <= x"06";
            when "01" & x"340" => data <= x"01";
            when "01" & x"341" => data <= x"a9";
            when "01" & x"342" => data <= x"06";
            when "01" & x"343" => data <= x"20";
            when "01" & x"344" => data <= x"15";
            when "01" & x"345" => data <= x"80";
            when "01" & x"346" => data <= x"a2";
            when "01" & x"347" => data <= x"0d";
            when "01" & x"348" => data <= x"bd";
            when "01" & x"349" => data <= x"49";
            when "01" & x"34a" => data <= x"99";
            when "01" & x"34b" => data <= x"9d";
            when "01" & x"34c" => data <= x"12";
            when "01" & x"34d" => data <= x"02";
            when "01" & x"34e" => data <= x"ca";
            when "01" & x"34f" => data <= x"10";
            when "01" & x"350" => data <= x"f7";
            when "01" & x"351" => data <= x"20";
            when "01" & x"352" => data <= x"28";
            when "01" & x"353" => data <= x"99";
            when "01" & x"354" => data <= x"84";
            when "01" & x"355" => data <= x"b1";
            when "01" & x"356" => data <= x"86";
            when "01" & x"357" => data <= x"b0";
            when "01" & x"358" => data <= x"a2";
            when "01" & x"359" => data <= x"07";
            when "01" & x"35a" => data <= x"a0";
            when "01" & x"35b" => data <= x"1b";
            when "01" & x"35c" => data <= x"b9";
            when "01" & x"35d" => data <= x"3c";
            when "01" & x"35e" => data <= x"99";
            when "01" & x"35f" => data <= x"91";
            when "01" & x"360" => data <= x"b0";
            when "01" & x"361" => data <= x"c8";
            when "01" & x"362" => data <= x"b9";
            when "01" & x"363" => data <= x"3c";
            when "01" & x"364" => data <= x"99";
            when "01" & x"365" => data <= x"91";
            when "01" & x"366" => data <= x"b0";
            when "01" & x"367" => data <= x"c8";
            when "01" & x"368" => data <= x"a5";
            when "01" & x"369" => data <= x"f4";
            when "01" & x"36a" => data <= x"91";
            when "01" & x"36b" => data <= x"b0";
            when "01" & x"36c" => data <= x"c8";
            when "01" & x"36d" => data <= x"ca";
            when "01" & x"36e" => data <= x"d0";
            when "01" & x"36f" => data <= x"ec";
            when "01" & x"370" => data <= x"86";
            when "01" & x"371" => data <= x"cf";
            when "01" & x"372" => data <= x"8c";
            when "01" & x"373" => data <= x"82";
            when "01" & x"374" => data <= x"10";
            when "01" & x"375" => data <= x"a2";
            when "01" & x"376" => data <= x"0f";
            when "01" & x"377" => data <= x"20";
            when "01" & x"378" => data <= x"2c";
            when "01" & x"379" => data <= x"99";
            when "01" & x"37a" => data <= x"20";
            when "01" & x"37b" => data <= x"9e";
            when "01" & x"37c" => data <= x"98";
            when "01" & x"37d" => data <= x"a0";
            when "01" & x"37e" => data <= x"d4";
            when "01" & x"37f" => data <= x"b1";
            when "01" & x"380" => data <= x"b0";
            when "01" & x"381" => data <= x"10";
            when "01" & x"382" => data <= x"2f";
            when "01" & x"383" => data <= x"a0";
            when "01" & x"384" => data <= x"d5";
            when "01" & x"385" => data <= x"b1";
            when "01" & x"386" => data <= x"b0";
            when "01" & x"387" => data <= x"30";
            when "01" & x"388" => data <= x"27";
            when "01" & x"389" => data <= x"20";
            when "01" & x"38a" => data <= x"8f";
            when "01" & x"38b" => data <= x"98";
            when "01" & x"38c" => data <= x"a0";
            when "01" & x"38d" => data <= x"00";
            when "01" & x"38e" => data <= x"b1";
            when "01" & x"38f" => data <= x"b0";
            when "01" & x"390" => data <= x"c0";
            when "01" & x"391" => data <= x"c0";
            when "01" & x"392" => data <= x"90";
            when "01" & x"393" => data <= x"05";
            when "01" & x"394" => data <= x"99";
            when "01" & x"395" => data <= x"00";
            when "01" & x"396" => data <= x"10";
            when "01" & x"397" => data <= x"b0";
            when "01" & x"398" => data <= x"03";
            when "01" & x"399" => data <= x"99";
            when "01" & x"39a" => data <= x"00";
            when "01" & x"39b" => data <= x"11";
            when "01" & x"39c" => data <= x"88";
            when "01" & x"39d" => data <= x"d0";
            when "01" & x"39e" => data <= x"ef";
            when "01" & x"39f" => data <= x"a9";
            when "01" & x"3a0" => data <= x"a0";
            when "01" & x"3a1" => data <= x"a8";
            when "01" & x"3a2" => data <= x"48";
            when "01" & x"3a3" => data <= x"a9";
            when "01" & x"3a4" => data <= x"3f";
            when "01" & x"3a5" => data <= x"20";
            when "01" & x"3a6" => data <= x"43";
            when "01" & x"3a7" => data <= x"91";
            when "01" & x"3a8" => data <= x"68";
            when "01" & x"3a9" => data <= x"99";
            when "01" & x"3aa" => data <= x"1d";
            when "01" & x"3ab" => data <= x"11";
            when "01" & x"3ac" => data <= x"e9";
            when "01" & x"3ad" => data <= x"1f";
            when "01" & x"3ae" => data <= x"d0";
            when "01" & x"3af" => data <= x"f1";
            when "01" & x"3b0" => data <= x"68";
            when "01" & x"3b1" => data <= x"60";
            when "01" & x"3b2" => data <= x"a9";
            when "01" & x"3b3" => data <= x"ff";
            when "01" & x"3b4" => data <= x"91";
            when "01" & x"3b5" => data <= x"b0";
            when "01" & x"3b6" => data <= x"8d";
            when "01" & x"3b7" => data <= x"d4";
            when "01" & x"3b8" => data <= x"10";
            when "01" & x"3b9" => data <= x"20";
            when "01" & x"3ba" => data <= x"8f";
            when "01" & x"3bb" => data <= x"98";
            when "01" & x"3bc" => data <= x"20";
            when "01" & x"3bd" => data <= x"24";
            when "01" & x"3be" => data <= x"99";
            when "01" & x"3bf" => data <= x"8a";
            when "01" & x"3c0" => data <= x"49";
            when "01" & x"3c1" => data <= x"ff";
            when "01" & x"3c2" => data <= x"8d";
            when "01" & x"3c3" => data <= x"d7";
            when "01" & x"3c4" => data <= x"10";
            when "01" & x"3c5" => data <= x"a9";
            when "01" & x"3c6" => data <= x"24";
            when "01" & x"3c7" => data <= x"8d";
            when "01" & x"3c8" => data <= x"ca";
            when "01" & x"3c9" => data <= x"10";
            when "01" & x"3ca" => data <= x"8d";
            when "01" & x"3cb" => data <= x"cc";
            when "01" & x"3cc" => data <= x"10";
            when "01" & x"3cd" => data <= x"a0";
            when "01" & x"3ce" => data <= x"00";
            when "01" & x"3cf" => data <= x"8c";
            when "01" & x"3d0" => data <= x"cb";
            when "01" & x"3d1" => data <= x"10";
            when "01" & x"3d2" => data <= x"8c";
            when "01" & x"3d3" => data <= x"cd";
            when "01" & x"3d4" => data <= x"10";
            when "01" & x"3d5" => data <= x"a0";
            when "01" & x"3d6" => data <= x"00";
            when "01" & x"3d7" => data <= x"8c";
            when "01" & x"3d8" => data <= x"c0";
            when "01" & x"3d9" => data <= x"10";
            when "01" & x"3da" => data <= x"8c";
            when "01" & x"3db" => data <= x"c9";
            when "01" & x"3dc" => data <= x"10";
            when "01" & x"3dd" => data <= x"88";
            when "01" & x"3de" => data <= x"8c";
            when "01" & x"3df" => data <= x"c8";
            when "01" & x"3e0" => data <= x"10";
            when "01" & x"3e1" => data <= x"8c";
            when "01" & x"3e2" => data <= x"c7";
            when "01" & x"3e3" => data <= x"10";
            when "01" & x"3e4" => data <= x"8c";
            when "01" & x"3e5" => data <= x"de";
            when "01" & x"3e6" => data <= x"10";
            when "01" & x"3e7" => data <= x"20";
            when "01" & x"3e8" => data <= x"37";
            when "01" & x"3e9" => data <= x"b1";
            when "01" & x"3ea" => data <= x"4c";
            when "01" & x"3eb" => data <= x"04";
            when "01" & x"3ec" => data <= x"94";
            when "01" & x"3ed" => data <= x"00";
            when "01" & x"3ee" => data <= x"00";
            when "01" & x"3ef" => data <= x"00";
            when "01" & x"3f0" => data <= x"00";
            when "01" & x"3f1" => data <= x"00";
            when "01" & x"3f2" => data <= x"00";
            when "01" & x"3f3" => data <= x"00";
            when "01" & x"3f4" => data <= x"00";
            when "01" & x"3f5" => data <= x"00";
            when "01" & x"3f6" => data <= x"00";
            when "01" & x"3f7" => data <= x"00";
            when "01" & x"3f8" => data <= x"00";
            when "01" & x"3f9" => data <= x"00";
            when "01" & x"3fa" => data <= x"00";
            when "01" & x"3fb" => data <= x"00";
            when "01" & x"3fc" => data <= x"00";
            when "01" & x"3fd" => data <= x"00";
            when "01" & x"3fe" => data <= x"00";
            when "01" & x"3ff" => data <= x"00";
            when "01" & x"400" => data <= x"00";
            when "01" & x"401" => data <= x"00";
            when "01" & x"402" => data <= x"00";
            when "01" & x"403" => data <= x"00";
            when "01" & x"404" => data <= x"68";
            when "01" & x"405" => data <= x"d0";
            when "01" & x"406" => data <= x"34";
            when "01" & x"407" => data <= x"20";
            when "01" & x"408" => data <= x"41";
            when "01" & x"409" => data <= x"af";
            when "01" & x"40a" => data <= x"a0";
            when "01" & x"40b" => data <= x"00";
            when "01" & x"40c" => data <= x"a2";
            when "01" & x"40d" => data <= x"00";
            when "01" & x"40e" => data <= x"ad";
            when "01" & x"40f" => data <= x"06";
            when "01" & x"410" => data <= x"0f";
            when "01" & x"411" => data <= x"20";
            when "01" & x"412" => data <= x"05";
            when "01" & x"413" => data <= x"82";
            when "01" & x"414" => data <= x"f0";
            when "01" & x"415" => data <= x"25";
            when "01" & x"416" => data <= x"48";
            when "01" & x"417" => data <= x"a2";
            when "01" & x"418" => data <= x"43";
            when "01" & x"419" => data <= x"a0";
            when "01" & x"41a" => data <= x"99";
            when "01" & x"41b" => data <= x"20";
            when "01" & x"41c" => data <= x"b8";
            when "01" & x"41d" => data <= x"86";
            when "01" & x"41e" => data <= x"20";
            when "01" & x"41f" => data <= x"fe";
            when "01" & x"420" => data <= x"80";
            when "01" & x"421" => data <= x"20";
            when "01" & x"422" => data <= x"96";
            when "01" & x"423" => data <= x"82";
            when "01" & x"424" => data <= x"68";
            when "01" & x"425" => data <= x"b0";
            when "01" & x"426" => data <= x"15";
            when "01" & x"427" => data <= x"20";
            when "01" & x"428" => data <= x"65";
            when "01" & x"429" => data <= x"80";
            when "01" & x"42a" => data <= x"46";
            when "01" & x"42b" => data <= x"69";
            when "01" & x"42c" => data <= x"6c";
            when "01" & x"42d" => data <= x"65";
            when "01" & x"42e" => data <= x"20";
            when "01" & x"42f" => data <= x"6e";
            when "01" & x"430" => data <= x"6f";
            when "01" & x"431" => data <= x"74";
            when "01" & x"432" => data <= x"20";
            when "01" & x"433" => data <= x"66";
            when "01" & x"434" => data <= x"6f";
            when "01" & x"435" => data <= x"75";
            when "01" & x"436" => data <= x"6e";
            when "01" & x"437" => data <= x"64";
            when "01" & x"438" => data <= x"0d";
            when "01" & x"439" => data <= x"0d";
            when "01" & x"43a" => data <= x"ea";
            when "01" & x"43b" => data <= x"60";
            when "01" & x"43c" => data <= x"c9";
            when "01" & x"43d" => data <= x"02";
            when "01" & x"43e" => data <= x"90";
            when "01" & x"43f" => data <= x"0e";
            when "01" & x"440" => data <= x"f0";
            when "01" & x"441" => data <= x"06";
            when "01" & x"442" => data <= x"a2";
            when "01" & x"443" => data <= x"41";
            when "01" & x"444" => data <= x"a0";
            when "01" & x"445" => data <= x"99";
            when "01" & x"446" => data <= x"d0";
            when "01" & x"447" => data <= x"0a";
            when "01" & x"448" => data <= x"a2";
            when "01" & x"449" => data <= x"43";
            when "01" & x"44a" => data <= x"a0";
            when "01" & x"44b" => data <= x"99";
            when "01" & x"44c" => data <= x"d0";
            when "01" & x"44d" => data <= x"04";
            when "01" & x"44e" => data <= x"a2";
            when "01" & x"44f" => data <= x"39";
            when "01" & x"450" => data <= x"a0";
            when "01" & x"451" => data <= x"99";
            when "01" & x"452" => data <= x"4c";
            when "01" & x"453" => data <= x"f7";
            when "01" & x"454" => data <= x"ff";
            when "01" & x"455" => data <= x"c9";
            when "01" & x"456" => data <= x"01";
            when "01" & x"457" => data <= x"d0";
            when "01" & x"458" => data <= x"07";
            when "01" & x"459" => data <= x"c0";
            when "01" & x"45a" => data <= x"17";
            when "01" & x"45b" => data <= x"b0";
            when "01" & x"45c" => data <= x"02";
            when "01" & x"45d" => data <= x"a0";
            when "01" & x"45e" => data <= x"17";
            when "01" & x"45f" => data <= x"60";
            when "01" & x"460" => data <= x"c9";
            when "01" & x"461" => data <= x"02";
            when "01" & x"462" => data <= x"d0";
            when "01" & x"463" => data <= x"1a";
            when "01" & x"464" => data <= x"48";
            when "01" & x"465" => data <= x"69";
            when "01" & x"466" => data <= x"12";
            when "01" & x"467" => data <= x"85";
            when "01" & x"468" => data <= x"b1";
            when "01" & x"469" => data <= x"9d";
            when "01" & x"46a" => data <= x"f0";
            when "01" & x"46b" => data <= x"0d";
            when "01" & x"46c" => data <= x"98";
            when "01" & x"46d" => data <= x"ea";
            when "01" & x"46e" => data <= x"48";
            when "01" & x"46f" => data <= x"a9";
            when "01" & x"470" => data <= x"00";
            when "01" & x"471" => data <= x"85";
            when "01" & x"472" => data <= x"b0";
            when "01" & x"473" => data <= x"a0";
            when "01" & x"474" => data <= x"d4";
            when "01" & x"475" => data <= x"91";
            when "01" & x"476" => data <= x"b0";
            when "01" & x"477" => data <= x"c8";
            when "01" & x"478" => data <= x"91";
            when "01" & x"479" => data <= x"b0";
            when "01" & x"47a" => data <= x"68";
            when "01" & x"47b" => data <= x"a8";
            when "01" & x"47c" => data <= x"68";
            when "01" & x"47d" => data <= x"60";
            when "01" & x"47e" => data <= x"c9";
            when "01" & x"47f" => data <= x"03";
            when "01" & x"480" => data <= x"d0";
            when "01" & x"481" => data <= x"19";
            when "01" & x"482" => data <= x"84";
            when "01" & x"483" => data <= x"b3";
            when "01" & x"484" => data <= x"20";
            when "01" & x"485" => data <= x"e1";
            when "01" & x"486" => data <= x"83";
            when "01" & x"487" => data <= x"4c";
            when "01" & x"488" => data <= x"8f";
            when "01" & x"489" => data <= x"a9";
            when "01" & x"48a" => data <= x"f4";
            when "01" & x"48b" => data <= x"ff";
            when "01" & x"48c" => data <= x"8a";
            when "01" & x"48d" => data <= x"30";
            when "01" & x"48e" => data <= x"09";
            when "01" & x"48f" => data <= x"c9";
            when "01" & x"490" => data <= x"32";
            when "01" & x"491" => data <= x"d0";
            when "01" & x"492" => data <= x"ea";
            when "01" & x"493" => data <= x"a9";
            when "01" & x"494" => data <= x"78";
            when "01" & x"495" => data <= x"20";
            when "01" & x"496" => data <= x"f4";
            when "01" & x"497" => data <= x"ff";
            when "01" & x"498" => data <= x"4c";
            when "01" & x"499" => data <= x"20";
            when "01" & x"49a" => data <= x"93";
            when "01" & x"49b" => data <= x"c9";
            when "01" & x"49c" => data <= x"04";
            when "01" & x"49d" => data <= x"d0";
            when "01" & x"49e" => data <= x"08";
            when "01" & x"49f" => data <= x"20";
            when "01" & x"4a0" => data <= x"e1";
            when "01" & x"4a1" => data <= x"83";
            when "01" & x"4a2" => data <= x"a2";
            when "01" & x"4a3" => data <= x"72";
            when "01" & x"4a4" => data <= x"4c";
            when "01" & x"4a5" => data <= x"71";
            when "01" & x"4a6" => data <= x"86";
            when "01" & x"4a7" => data <= x"c9";
            when "01" & x"4a8" => data <= x"09";
            when "01" & x"4a9" => data <= x"d0";
            when "01" & x"4aa" => data <= x"12";
            when "01" & x"4ab" => data <= x"20";
            when "01" & x"4ac" => data <= x"e1";
            when "01" & x"4ad" => data <= x"83";
            when "01" & x"4ae" => data <= x"4c";
            when "01" & x"4af" => data <= x"cc";
            when "01" & x"4b0" => data <= x"b3";
            when "01" & x"4b1" => data <= x"a0";
            when "01" & x"4b2" => data <= x"c9";
            when "01" & x"4b3" => data <= x"0d";
            when "01" & x"4b4" => data <= x"d0";
            when "01" & x"4b5" => data <= x"ee";
            when "01" & x"4b6" => data <= x"98";
            when "01" & x"4b7" => data <= x"e8";
            when "01" & x"4b8" => data <= x"a0";
            when "01" & x"4b9" => data <= x"02";
            when "01" & x"4ba" => data <= x"4c";
            when "01" & x"4bb" => data <= x"cb";
            when "01" & x"4bc" => data <= x"99";
            when "01" & x"4bd" => data <= x"c9";
            when "01" & x"4be" => data <= x"0a";
            when "01" & x"4bf" => data <= x"d0";
            when "01" & x"4c0" => data <= x"29";
            when "01" & x"4c1" => data <= x"20";
            when "01" & x"4c2" => data <= x"e1";
            when "01" & x"4c3" => data <= x"83";
            when "01" & x"4c4" => data <= x"20";
            when "01" & x"4c5" => data <= x"9e";
            when "01" & x"4c6" => data <= x"98";
            when "01" & x"4c7" => data <= x"a0";
            when "01" & x"4c8" => data <= x"d5";
            when "01" & x"4c9" => data <= x"b1";
            when "01" & x"4ca" => data <= x"b0";
            when "01" & x"4cb" => data <= x"10";
            when "01" & x"4cc" => data <= x"1c";
            when "01" & x"4cd" => data <= x"a0";
            when "01" & x"4ce" => data <= x"00";
            when "01" & x"4cf" => data <= x"c0";
            when "01" & x"4d0" => data <= x"c0";
            when "01" & x"4d1" => data <= x"90";
            when "01" & x"4d2" => data <= x"05";
            when "01" & x"4d3" => data <= x"b9";
            when "01" & x"4d4" => data <= x"00";
            when "01" & x"4d5" => data <= x"10";
            when "01" & x"4d6" => data <= x"b0";
            when "01" & x"4d7" => data <= x"03";
            when "01" & x"4d8" => data <= x"b9";
            when "01" & x"4d9" => data <= x"00";
            when "01" & x"4da" => data <= x"11";
            when "01" & x"4db" => data <= x"91";
            when "01" & x"4dc" => data <= x"b0";
            when "01" & x"4dd" => data <= x"88";
            when "01" & x"4de" => data <= x"d0";
            when "01" & x"4df" => data <= x"ef";
            when "01" & x"4e0" => data <= x"20";
            when "01" & x"4e1" => data <= x"f2";
            when "01" & x"4e2" => data <= x"8f";
            when "01" & x"4e3" => data <= x"a0";
            when "01" & x"4e4" => data <= x"d5";
            when "01" & x"4e5" => data <= x"a9";
            when "01" & x"4e6" => data <= x"00";
            when "01" & x"4e7" => data <= x"91";
            when "01" & x"4e8" => data <= x"b0";
            when "01" & x"4e9" => data <= x"60";
            when "01" & x"4ea" => data <= x"c9";
            when "01" & x"4eb" => data <= x"08";
            when "01" & x"4ec" => data <= x"d0";
            when "01" & x"4ed" => data <= x"15";
            when "01" & x"4ee" => data <= x"20";
            when "01" & x"4ef" => data <= x"11";
            when "01" & x"4f0" => data <= x"84";
            when "01" & x"4f1" => data <= x"a4";
            when "01" & x"4f2" => data <= x"f0";
            when "01" & x"4f3" => data <= x"84";
            when "01" & x"4f4" => data <= x"b0";
            when "01" & x"4f5" => data <= x"a4";
            when "01" & x"4f6" => data <= x"f1";
            when "01" & x"4f7" => data <= x"84";
            when "01" & x"4f8" => data <= x"b1";
            when "01" & x"4f9" => data <= x"a4";
            when "01" & x"4fa" => data <= x"ef";
            when "01" & x"4fb" => data <= x"c0";
            when "01" & x"4fc" => data <= x"7f";
            when "01" & x"4fd" => data <= x"d0";
            when "01" & x"4fe" => data <= x"4c";
            when "01" & x"4ff" => data <= x"4c";
            when "01" & x"500" => data <= x"46";
            when "01" & x"501" => data <= x"be";
            when "01" & x"502" => data <= x"00";
            when "01" & x"503" => data <= x"4c";
            when "01" & x"504" => data <= x"f6";
            when "01" & x"505" => data <= x"a0";
            when "01" & x"506" => data <= x"00";
            when "01" & x"507" => data <= x"00";
            when "01" & x"508" => data <= x"00";
            when "01" & x"509" => data <= x"00";
            when "01" & x"50a" => data <= x"00";
            when "01" & x"50b" => data <= x"00";
            when "01" & x"50c" => data <= x"00";
            when "01" & x"50d" => data <= x"00";
            when "01" & x"50e" => data <= x"00";
            when "01" & x"50f" => data <= x"00";
            when "01" & x"510" => data <= x"00";
            when "01" & x"511" => data <= x"00";
            when "01" & x"512" => data <= x"00";
            when "01" & x"513" => data <= x"00";
            when "01" & x"514" => data <= x"00";
            when "01" & x"515" => data <= x"00";
            when "01" & x"516" => data <= x"00";
            when "01" & x"517" => data <= x"00";
            when "01" & x"518" => data <= x"00";
            when "01" & x"519" => data <= x"00";
            when "01" & x"51a" => data <= x"00";
            when "01" & x"51b" => data <= x"00";
            when "01" & x"51c" => data <= x"00";
            when "01" & x"51d" => data <= x"00";
            when "01" & x"51e" => data <= x"00";
            when "01" & x"51f" => data <= x"00";
            when "01" & x"520" => data <= x"00";
            when "01" & x"521" => data <= x"00";
            when "01" & x"522" => data <= x"00";
            when "01" & x"523" => data <= x"00";
            when "01" & x"524" => data <= x"00";
            when "01" & x"525" => data <= x"00";
            when "01" & x"526" => data <= x"00";
            when "01" & x"527" => data <= x"00";
            when "01" & x"528" => data <= x"00";
            when "01" & x"529" => data <= x"00";
            when "01" & x"52a" => data <= x"00";
            when "01" & x"52b" => data <= x"00";
            when "01" & x"52c" => data <= x"00";
            when "01" & x"52d" => data <= x"00";
            when "01" & x"52e" => data <= x"00";
            when "01" & x"52f" => data <= x"00";
            when "01" & x"530" => data <= x"00";
            when "01" & x"531" => data <= x"00";
            when "01" & x"532" => data <= x"00";
            when "01" & x"533" => data <= x"00";
            when "01" & x"534" => data <= x"00";
            when "01" & x"535" => data <= x"00";
            when "01" & x"536" => data <= x"00";
            when "01" & x"537" => data <= x"00";
            when "01" & x"538" => data <= x"00";
            when "01" & x"539" => data <= x"00";
            when "01" & x"53a" => data <= x"00";
            when "01" & x"53b" => data <= x"00";
            when "01" & x"53c" => data <= x"00";
            when "01" & x"53d" => data <= x"00";
            when "01" & x"53e" => data <= x"00";
            when "01" & x"53f" => data <= x"00";
            when "01" & x"540" => data <= x"00";
            when "01" & x"541" => data <= x"00";
            when "01" & x"542" => data <= x"00";
            when "01" & x"543" => data <= x"00";
            when "01" & x"544" => data <= x"00";
            when "01" & x"545" => data <= x"00";
            when "01" & x"546" => data <= x"00";
            when "01" & x"547" => data <= x"00";
            when "01" & x"548" => data <= x"00";
            when "01" & x"549" => data <= x"00";
            when "01" & x"54a" => data <= x"00";
            when "01" & x"54b" => data <= x"c0";
            when "01" & x"54c" => data <= x"7d";
            when "01" & x"54d" => data <= x"90";
            when "01" & x"54e" => data <= x"2b";
            when "01" & x"54f" => data <= x"20";
            when "01" & x"550" => data <= x"4d";
            when "01" & x"551" => data <= x"83";
            when "01" & x"552" => data <= x"20";
            when "01" & x"553" => data <= x"47";
            when "01" & x"554" => data <= x"83";
            when "01" & x"555" => data <= x"c0";
            when "01" & x"556" => data <= x"7e";
            when "01" & x"557" => data <= x"f0";
            when "01" & x"558" => data <= x"09";
            when "01" & x"559" => data <= x"a0";
            when "01" & x"55a" => data <= x"00";
            when "01" & x"55b" => data <= x"ad";
            when "01" & x"55c" => data <= x"04";
            when "01" & x"55d" => data <= x"0f";
            when "01" & x"55e" => data <= x"91";
            when "01" & x"55f" => data <= x"b0";
            when "01" & x"560" => data <= x"98";
            when "01" & x"561" => data <= x"60";
            when "01" & x"562" => data <= x"a9";
            when "01" & x"563" => data <= x"00";
            when "01" & x"564" => data <= x"a8";
            when "01" & x"565" => data <= x"91";
            when "01" & x"566" => data <= x"b0";
            when "01" & x"567" => data <= x"c8";
            when "01" & x"568" => data <= x"ad";
            when "01" & x"569" => data <= x"07";
            when "01" & x"56a" => data <= x"0f";
            when "01" & x"56b" => data <= x"91";
            when "01" & x"56c" => data <= x"b0";
            when "01" & x"56d" => data <= x"c8";
            when "01" & x"56e" => data <= x"ad";
            when "01" & x"56f" => data <= x"06";
            when "01" & x"570" => data <= x"0f";
            when "01" & x"571" => data <= x"29";
            when "01" & x"572" => data <= x"03";
            when "01" & x"573" => data <= x"91";
            when "01" & x"574" => data <= x"b0";
            when "01" & x"575" => data <= x"c8";
            when "01" & x"576" => data <= x"a9";
            when "01" & x"577" => data <= x"00";
            when "01" & x"578" => data <= x"91";
            when "01" & x"579" => data <= x"b0";
            when "01" & x"57a" => data <= x"60";
            when "01" & x"57b" => data <= x"20";
            when "01" & x"57c" => data <= x"11";
            when "01" & x"57d" => data <= x"84";
            when "01" & x"57e" => data <= x"48";
            when "01" & x"57f" => data <= x"20";
            when "01" & x"580" => data <= x"62";
            when "01" & x"581" => data <= x"82";
            when "01" & x"582" => data <= x"86";
            when "01" & x"583" => data <= x"b0";
            when "01" & x"584" => data <= x"8e";
            when "01" & x"585" => data <= x"dc";
            when "01" & x"586" => data <= x"10";
            when "01" & x"587" => data <= x"84";
            when "01" & x"588" => data <= x"b1";
            when "01" & x"589" => data <= x"8c";
            when "01" & x"58a" => data <= x"dd";
            when "01" & x"58b" => data <= x"10";
            when "01" & x"58c" => data <= x"a2";
            when "01" & x"58d" => data <= x"00";
            when "01" & x"58e" => data <= x"a0";
            when "01" & x"58f" => data <= x"00";
            when "01" & x"590" => data <= x"20";
            when "01" & x"591" => data <= x"ea";
            when "01" & x"592" => data <= x"80";
            when "01" & x"593" => data <= x"20";
            when "01" & x"594" => data <= x"da";
            when "01" & x"595" => data <= x"80";
            when "01" & x"596" => data <= x"c0";
            when "01" & x"597" => data <= x"12";
            when "01" & x"598" => data <= x"d0";
            when "01" & x"599" => data <= x"f9";
            when "01" & x"59a" => data <= x"68";
            when "01" & x"59b" => data <= x"aa";
            when "01" & x"59c" => data <= x"e8";
            when "01" & x"59d" => data <= x"e0";
            when "01" & x"59e" => data <= x"08";
            when "01" & x"59f" => data <= x"b0";
            when "01" & x"5a0" => data <= x"08";
            when "01" & x"5a1" => data <= x"bd";
            when "01" & x"5a2" => data <= x"8c";
            when "01" & x"5a3" => data <= x"99";
            when "01" & x"5a4" => data <= x"48";
            when "01" & x"5a5" => data <= x"bd";
            when "01" & x"5a6" => data <= x"84";
            when "01" & x"5a7" => data <= x"99";
            when "01" & x"5a8" => data <= x"48";
            when "01" & x"5a9" => data <= x"60";
            when "01" & x"5aa" => data <= x"c9";
            when "01" & x"5ab" => data <= x"09";
            when "01" & x"5ac" => data <= x"b0";
            when "01" & x"5ad" => data <= x"fb";
            when "01" & x"5ae" => data <= x"86";
            when "01" & x"5af" => data <= x"b5";
            when "01" & x"5b0" => data <= x"aa";
            when "01" & x"5b1" => data <= x"bd";
            when "01" & x"5b2" => data <= x"75";
            when "01" & x"5b3" => data <= x"99";
            when "01" & x"5b4" => data <= x"48";
            when "01" & x"5b5" => data <= x"bd";
            when "01" & x"5b6" => data <= x"6c";
            when "01" & x"5b7" => data <= x"99";
            when "01" & x"5b8" => data <= x"48";
            when "01" & x"5b9" => data <= x"8a";
            when "01" & x"5ba" => data <= x"a6";
            when "01" & x"5bb" => data <= x"b5";
            when "01" & x"5bc" => data <= x"60";
            when "01" & x"5bd" => data <= x"a9";
            when "01" & x"5be" => data <= x"ff";
            when "01" & x"5bf" => data <= x"95";
            when "01" & x"5c0" => data <= x"02";
            when "01" & x"5c1" => data <= x"95";
            when "01" & x"5c2" => data <= x"03";
            when "01" & x"5c3" => data <= x"ad";
            when "01" & x"5c4" => data <= x"da";
            when "01" & x"5c5" => data <= x"10";
            when "01" & x"5c6" => data <= x"95";
            when "01" & x"5c7" => data <= x"00";
            when "01" & x"5c8" => data <= x"ad";
            when "01" & x"5c9" => data <= x"db";
            when "01" & x"5ca" => data <= x"10";
            when "01" & x"5cb" => data <= x"95";
            when "01" & x"5cc" => data <= x"01";
            when "01" & x"5cd" => data <= x"a9";
            when "01" & x"5ce" => data <= x"00";
            when "01" & x"5cf" => data <= x"60";
            when "01" & x"5d0" => data <= x"c9";
            when "01" & x"5d1" => data <= x"09";
            when "01" & x"5d2" => data <= x"b0";
            when "01" & x"5d3" => data <= x"fb";
            when "01" & x"5d4" => data <= x"20";
            when "01" & x"5d5" => data <= x"e1";
            when "01" & x"5d6" => data <= x"83";
            when "01" & x"5d7" => data <= x"8e";
            when "01" & x"5d8" => data <= x"7d";
            when "01" & x"5d9" => data <= x"10";
            when "01" & x"5da" => data <= x"8c";
            when "01" & x"5db" => data <= x"7e";
            when "01" & x"5dc" => data <= x"10";
            when "01" & x"5dd" => data <= x"a8";
            when "01" & x"5de" => data <= x"ba";
            when "01" & x"5df" => data <= x"a9";
            when "01" & x"5e0" => data <= x"00";
            when "01" & x"5e1" => data <= x"4c";
            when "01" & x"5e2" => data <= x"d8";
            when "01" & x"5e3" => data <= x"a0";
            when "01" & x"5e4" => data <= x"b9";
            when "01" & x"5e5" => data <= x"ab";
            when "01" & x"5e6" => data <= x"99";
            when "01" & x"5e7" => data <= x"8d";
            when "01" & x"5e8" => data <= x"d8";
            when "01" & x"5e9" => data <= x"10";
            when "01" & x"5ea" => data <= x"b9";
            when "01" & x"5eb" => data <= x"b4";
            when "01" & x"5ec" => data <= x"99";
            when "01" & x"5ed" => data <= x"8d";
            when "01" & x"5ee" => data <= x"d9";
            when "01" & x"5ef" => data <= x"10";
            when "01" & x"5f0" => data <= x"b9";
            when "01" & x"5f1" => data <= x"bd";
            when "01" & x"5f2" => data <= x"99";
            when "01" & x"5f3" => data <= x"4a";
            when "01" & x"5f4" => data <= x"08";
            when "01" & x"5f5" => data <= x"4a";
            when "01" & x"5f6" => data <= x"08";
            when "01" & x"5f7" => data <= x"8d";
            when "01" & x"5f8" => data <= x"7f";
            when "01" & x"5f9" => data <= x"10";
            when "01" & x"5fa" => data <= x"20";
            when "01" & x"5fb" => data <= x"56";
            when "01" & x"5fc" => data <= x"97";
            when "01" & x"5fd" => data <= x"a0";
            when "01" & x"5fe" => data <= x"0c";
            when "01" & x"5ff" => data <= x"b1";
            when "01" & x"600" => data <= x"b4";
            when "01" & x"601" => data <= x"99";
            when "01" & x"602" => data <= x"60";
            when "01" & x"603" => data <= x"10";
            when "01" & x"604" => data <= x"88";
            when "01" & x"605" => data <= x"10";
            when "01" & x"606" => data <= x"f8";
            when "01" & x"607" => data <= x"ad";
            when "01" & x"608" => data <= x"63";
            when "01" & x"609" => data <= x"10";
            when "01" & x"60a" => data <= x"2d";
            when "01" & x"60b" => data <= x"64";
            when "01" & x"60c" => data <= x"10";
            when "01" & x"60d" => data <= x"0d";
            when "01" & x"60e" => data <= x"d7";
            when "01" & x"60f" => data <= x"10";
            when "01" & x"610" => data <= x"18";
            when "01" & x"611" => data <= x"69";
            when "01" & x"612" => data <= x"01";
            when "01" & x"613" => data <= x"4c";
            when "01" & x"614" => data <= x"eb";
            when "01" & x"615" => data <= x"a0";
            when "01" & x"616" => data <= x"ea";
            when "01" & x"617" => data <= x"8d";
            when "01" & x"618" => data <= x"81";
            when "01" & x"619" => data <= x"10";
            when "01" & x"61a" => data <= x"ad";
            when "01" & x"61b" => data <= x"7f";
            when "01" & x"61c" => data <= x"10";
            when "01" & x"61d" => data <= x"b0";
            when "01" & x"61e" => data <= x"07";
            when "01" & x"61f" => data <= x"a2";
            when "01" & x"620" => data <= x"61";
            when "01" & x"621" => data <= x"a0";
            when "01" & x"622" => data <= x"10";
            when "01" & x"623" => data <= x"20";
            when "01" & x"624" => data <= x"06";
            when "01" & x"625" => data <= x"04";
            when "01" & x"626" => data <= x"28";
            when "01" & x"627" => data <= x"b0";
            when "01" & x"628" => data <= x"04";
            when "01" & x"629" => data <= x"28";
            when "01" & x"62a" => data <= x"6c";
            when "01" & x"62b" => data <= x"d8";
            when "01" & x"62c" => data <= x"10";
            when "01" & x"62d" => data <= x"a2";
            when "01" & x"62e" => data <= x"03";
            when "01" & x"62f" => data <= x"bd";
            when "01" & x"630" => data <= x"69";
            when "01" & x"631" => data <= x"10";
            when "01" & x"632" => data <= x"95";
            when "01" & x"633" => data <= x"b6";
            when "01" & x"634" => data <= x"ca";
            when "01" & x"635" => data <= x"10";
            when "01" & x"636" => data <= x"f8";
            when "01" & x"637" => data <= x"a2";
            when "01" & x"638" => data <= x"b6";
            when "01" & x"639" => data <= x"ac";
            when "01" & x"63a" => data <= x"60";
            when "01" & x"63b" => data <= x"10";
            when "01" & x"63c" => data <= x"a9";
            when "01" & x"63d" => data <= x"00";
            when "01" & x"63e" => data <= x"28";
            when "01" & x"63f" => data <= x"b0";
            when "01" & x"640" => data <= x"03";
            when "01" & x"641" => data <= x"20";
            when "01" & x"642" => data <= x"a7";
            when "01" & x"643" => data <= x"92";
            when "01" & x"644" => data <= x"20";
            when "01" & x"645" => data <= x"2e";
            when "01" & x"646" => data <= x"90";
            when "01" & x"647" => data <= x"a2";
            when "01" & x"648" => data <= x"03";
            when "01" & x"649" => data <= x"b5";
            when "01" & x"64a" => data <= x"b6";
            when "01" & x"64b" => data <= x"9d";
            when "01" & x"64c" => data <= x"69";
            when "01" & x"64d" => data <= x"10";
            when "01" & x"64e" => data <= x"ca";
            when "01" & x"64f" => data <= x"10";
            when "01" & x"650" => data <= x"f8";
            when "01" & x"651" => data <= x"20";
            when "01" & x"652" => data <= x"48";
            when "01" & x"653" => data <= x"97";
            when "01" & x"654" => data <= x"30";
            when "01" & x"655" => data <= x"0d";
            when "01" & x"656" => data <= x"ac";
            when "01" & x"657" => data <= x"60";
            when "01" & x"658" => data <= x"10";
            when "01" & x"659" => data <= x"20";
            when "01" & x"65a" => data <= x"2a";
            when "01" & x"65b" => data <= x"96";
            when "01" & x"65c" => data <= x"b0";
            when "01" & x"65d" => data <= x"0d";
            when "01" & x"65e" => data <= x"a2";
            when "01" & x"65f" => data <= x"09";
            when "01" & x"660" => data <= x"20";
            when "01" & x"661" => data <= x"3c";
            when "01" & x"662" => data <= x"97";
            when "01" & x"663" => data <= x"a2";
            when "01" & x"664" => data <= x"05";
            when "01" & x"665" => data <= x"20";
            when "01" & x"666" => data <= x"3c";
            when "01" & x"667" => data <= x"97";
            when "01" & x"668" => data <= x"d0";
            when "01" & x"669" => data <= x"ec";
            when "01" & x"66a" => data <= x"18";
            when "01" & x"66b" => data <= x"08";
            when "01" & x"66c" => data <= x"20";
            when "01" & x"66d" => data <= x"48";
            when "01" & x"66e" => data <= x"97";
            when "01" & x"66f" => data <= x"a2";
            when "01" & x"670" => data <= x"05";
            when "01" & x"671" => data <= x"20";
            when "01" & x"672" => data <= x"3c";
            when "01" & x"673" => data <= x"97";
            when "01" & x"674" => data <= x"a0";
            when "01" & x"675" => data <= x"0c";
            when "01" & x"676" => data <= x"20";
            when "01" & x"677" => data <= x"56";
            when "01" & x"678" => data <= x"97";
            when "01" & x"679" => data <= x"b9";
            when "01" & x"67a" => data <= x"60";
            when "01" & x"67b" => data <= x"10";
            when "01" & x"67c" => data <= x"91";
            when "01" & x"67d" => data <= x"b4";
            when "01" & x"67e" => data <= x"88";
            when "01" & x"67f" => data <= x"10";
            when "01" & x"680" => data <= x"f8";
            when "01" & x"681" => data <= x"28";
            when "01" & x"682" => data <= x"60";
            when "01" & x"683" => data <= x"20";
            when "01" & x"684" => data <= x"4d";
            when "01" & x"685" => data <= x"83";
            when "01" & x"686" => data <= x"20";
            when "01" & x"687" => data <= x"41";
            when "01" & x"688" => data <= x"af";
            when "01" & x"689" => data <= x"a9";
            when "01" & x"68a" => data <= x"95";
            when "01" & x"68b" => data <= x"8d";
            when "01" & x"68c" => data <= x"d8";
            when "01" & x"68d" => data <= x"10";
            when "01" & x"68e" => data <= x"a9";
            when "01" & x"68f" => data <= x"96";
            when "01" & x"690" => data <= x"8d";
            when "01" & x"691" => data <= x"d9";
            when "01" & x"692" => data <= x"10";
            when "01" & x"693" => data <= x"d0";
            when "01" & x"694" => data <= x"bc";
            when "01" & x"695" => data <= x"ac";
            when "01" & x"696" => data <= x"69";
            when "01" & x"697" => data <= x"10";
            when "01" & x"698" => data <= x"cc";
            when "01" & x"699" => data <= x"05";
            when "01" & x"69a" => data <= x"0f";
            when "01" & x"69b" => data <= x"b0";
            when "01" & x"69c" => data <= x"28";
            when "01" & x"69d" => data <= x"b9";
            when "01" & x"69e" => data <= x"0f";
            when "01" & x"69f" => data <= x"0e";
            when "01" & x"6a0" => data <= x"20";
            when "01" & x"6a1" => data <= x"ee";
            when "01" & x"6a2" => data <= x"82";
            when "01" & x"6a3" => data <= x"45";
            when "01" & x"6a4" => data <= x"ce";
            when "01" & x"6a5" => data <= x"b0";
            when "01" & x"6a6" => data <= x"02";
            when "01" & x"6a7" => data <= x"29";
            when "01" & x"6a8" => data <= x"df";
            when "01" & x"6a9" => data <= x"29";
            when "01" & x"6aa" => data <= x"7f";
            when "01" & x"6ab" => data <= x"f0";
            when "01" & x"6ac" => data <= x"05";
            when "01" & x"6ad" => data <= x"20";
            when "01" & x"6ae" => data <= x"10";
            when "01" & x"6af" => data <= x"82";
            when "01" & x"6b0" => data <= x"d0";
            when "01" & x"6b1" => data <= x"e6";
            when "01" & x"6b2" => data <= x"a9";
            when "01" & x"6b3" => data <= x"07";
            when "01" & x"6b4" => data <= x"20";
            when "01" & x"6b5" => data <= x"6a";
            when "01" & x"6b6" => data <= x"97";
            when "01" & x"6b7" => data <= x"85";
            when "01" & x"6b8" => data <= x"b0";
            when "01" & x"6b9" => data <= x"b9";
            when "01" & x"6ba" => data <= x"08";
            when "01" & x"6bb" => data <= x"0e";
            when "01" & x"6bc" => data <= x"20";
            when "01" & x"6bd" => data <= x"6a";
            when "01" & x"6be" => data <= x"97";
            when "01" & x"6bf" => data <= x"c8";
            when "01" & x"6c0" => data <= x"c6";
            when "01" & x"6c1" => data <= x"b0";
            when "01" & x"6c2" => data <= x"d0";
            when "01" & x"6c3" => data <= x"f5";
            when "01" & x"6c4" => data <= x"18";
            when "01" & x"6c5" => data <= x"8c";
            when "01" & x"6c6" => data <= x"69";
            when "01" & x"6c7" => data <= x"10";
            when "01" & x"6c8" => data <= x"ad";
            when "01" & x"6c9" => data <= x"04";
            when "01" & x"6ca" => data <= x"0f";
            when "01" & x"6cb" => data <= x"8d";
            when "01" & x"6cc" => data <= x"60";
            when "01" & x"6cd" => data <= x"10";
            when "01" & x"6ce" => data <= x"60";
            when "01" & x"6cf" => data <= x"20";
            when "01" & x"6d0" => data <= x"4d";
            when "01" & x"6d1" => data <= x"83";
            when "01" & x"6d2" => data <= x"20";
            when "01" & x"6d3" => data <= x"41";
            when "01" & x"6d4" => data <= x"af";
            when "01" & x"6d5" => data <= x"a9";
            when "01" & x"6d6" => data <= x"0c";
            when "01" & x"6d7" => data <= x"20";
            when "01" & x"6d8" => data <= x"6a";
            when "01" & x"6d9" => data <= x"97";
            when "01" & x"6da" => data <= x"a0";
            when "01" & x"6db" => data <= x"00";
            when "01" & x"6dc" => data <= x"b9";
            when "01" & x"6dd" => data <= x"00";
            when "01" & x"6de" => data <= x"0e";
            when "01" & x"6df" => data <= x"20";
            when "01" & x"6e0" => data <= x"6a";
            when "01" & x"6e1" => data <= x"97";
            when "01" & x"6e2" => data <= x"c8";
            when "01" & x"6e3" => data <= x"c0";
            when "01" & x"6e4" => data <= x"08";
            when "01" & x"6e5" => data <= x"d0";
            when "01" & x"6e6" => data <= x"f5";
            when "01" & x"6e7" => data <= x"b9";
            when "01" & x"6e8" => data <= x"f8";
            when "01" & x"6e9" => data <= x"0e";
            when "01" & x"6ea" => data <= x"20";
            when "01" & x"6eb" => data <= x"6a";
            when "01" & x"6ec" => data <= x"97";
            when "01" & x"6ed" => data <= x"c8";
            when "01" & x"6ee" => data <= x"c0";
            when "01" & x"6ef" => data <= x"0c";
            when "01" & x"6f0" => data <= x"d0";
            when "01" & x"6f1" => data <= x"f5";
            when "01" & x"6f2" => data <= x"ad";
            when "01" & x"6f3" => data <= x"06";
            when "01" & x"6f4" => data <= x"0f";
            when "01" & x"6f5" => data <= x"20";
            when "01" & x"6f6" => data <= x"05";
            when "01" & x"6f7" => data <= x"82";
            when "01" & x"6f8" => data <= x"20";
            when "01" & x"6f9" => data <= x"6a";
            when "01" & x"6fa" => data <= x"97";
            when "01" & x"6fb" => data <= x"a5";
            when "01" & x"6fc" => data <= x"cf";
            when "01" & x"6fd" => data <= x"4c";
            when "01" & x"6fe" => data <= x"6a";
            when "01" & x"6ff" => data <= x"97";
            when "01" & x"700" => data <= x"20";
            when "01" & x"701" => data <= x"61";
            when "01" & x"702" => data <= x"97";
            when "01" & x"703" => data <= x"ad";
            when "01" & x"704" => data <= x"cb";
            when "01" & x"705" => data <= x"10";
            when "01" & x"706" => data <= x"09";
            when "01" & x"707" => data <= x"30";
            when "01" & x"708" => data <= x"20";
            when "01" & x"709" => data <= x"6a";
            when "01" & x"70a" => data <= x"97";
            when "01" & x"70b" => data <= x"20";
            when "01" & x"70c" => data <= x"61";
            when "01" & x"70d" => data <= x"97";
            when "01" & x"70e" => data <= x"ad";
            when "01" & x"70f" => data <= x"ca";
            when "01" & x"710" => data <= x"10";
            when "01" & x"711" => data <= x"4c";
            when "01" & x"712" => data <= x"6a";
            when "01" & x"713" => data <= x"97";
            when "01" & x"714" => data <= x"20";
            when "01" & x"715" => data <= x"61";
            when "01" & x"716" => data <= x"97";
            when "01" & x"717" => data <= x"ad";
            when "01" & x"718" => data <= x"cd";
            when "01" & x"719" => data <= x"10";
            when "01" & x"71a" => data <= x"09";
            when "01" & x"71b" => data <= x"30";
            when "01" & x"71c" => data <= x"20";
            when "01" & x"71d" => data <= x"6a";
            when "01" & x"71e" => data <= x"97";
            when "01" & x"71f" => data <= x"20";
            when "01" & x"720" => data <= x"61";
            when "01" & x"721" => data <= x"97";
            when "01" & x"722" => data <= x"ad";
            when "01" & x"723" => data <= x"cc";
            when "01" & x"724" => data <= x"10";
            when "01" & x"725" => data <= x"4c";
            when "01" & x"726" => data <= x"6a";
            when "01" & x"727" => data <= x"97";
            when "01" & x"728" => data <= x"48";
            when "01" & x"729" => data <= x"ad";
            when "01" & x"72a" => data <= x"61";
            when "01" & x"72b" => data <= x"10";
            when "01" & x"72c" => data <= x"85";
            when "01" & x"72d" => data <= x"b8";
            when "01" & x"72e" => data <= x"ad";
            when "01" & x"72f" => data <= x"62";
            when "01" & x"730" => data <= x"10";
            when "01" & x"731" => data <= x"85";
            when "01" & x"732" => data <= x"b9";
            when "01" & x"733" => data <= x"a2";
            when "01" & x"734" => data <= x"00";
            when "01" & x"735" => data <= x"68";
            when "01" & x"736" => data <= x"60";
            when "01" & x"737" => data <= x"20";
            when "01" & x"738" => data <= x"e1";
            when "01" & x"739" => data <= x"83";
            when "01" & x"73a" => data <= x"a2";
            when "01" & x"73b" => data <= x"01";
            when "01" & x"73c" => data <= x"a0";
            when "01" & x"73d" => data <= x"04";
            when "01" & x"73e" => data <= x"fe";
            when "01" & x"73f" => data <= x"60";
            when "01" & x"740" => data <= x"10";
            when "01" & x"741" => data <= x"d0";
            when "01" & x"742" => data <= x"04";
            when "01" & x"743" => data <= x"e8";
            when "01" & x"744" => data <= x"88";
            when "01" & x"745" => data <= x"d0";
            when "01" & x"746" => data <= x"f7";
            when "01" & x"747" => data <= x"60";
            when "01" & x"748" => data <= x"a2";
            when "01" & x"749" => data <= x"03";
            when "01" & x"74a" => data <= x"a9";
            when "01" & x"74b" => data <= x"ff";
            when "01" & x"74c" => data <= x"5d";
            when "01" & x"74d" => data <= x"65";
            when "01" & x"74e" => data <= x"10";
            when "01" & x"74f" => data <= x"9d";
            when "01" & x"750" => data <= x"65";
            when "01" & x"751" => data <= x"10";
            when "01" & x"752" => data <= x"ca";
            when "01" & x"753" => data <= x"10";
            when "01" & x"754" => data <= x"f5";
            when "01" & x"755" => data <= x"60";
            when "01" & x"756" => data <= x"ad";
            when "01" & x"757" => data <= x"7d";
            when "01" & x"758" => data <= x"10";
            when "01" & x"759" => data <= x"85";
            when "01" & x"75a" => data <= x"b4";
            when "01" & x"75b" => data <= x"ad";
            when "01" & x"75c" => data <= x"7e";
            when "01" & x"75d" => data <= x"10";
            when "01" & x"75e" => data <= x"85";
            when "01" & x"75f" => data <= x"b5";
            when "01" & x"760" => data <= x"60";
            when "01" & x"761" => data <= x"a9";
            when "01" & x"762" => data <= x"01";
            when "01" & x"763" => data <= x"d0";
            when "01" & x"764" => data <= x"05";
            when "01" & x"765" => data <= x"20";
            when "01" & x"766" => data <= x"c1";
            when "01" & x"767" => data <= x"90";
            when "01" & x"768" => data <= x"b0";
            when "01" & x"769" => data <= x"f6";
            when "01" & x"76a" => data <= x"2c";
            when "01" & x"76b" => data <= x"81";
            when "01" & x"76c" => data <= x"10";
            when "01" & x"76d" => data <= x"10";
            when "01" & x"76e" => data <= x"06";
            when "01" & x"76f" => data <= x"8d";
            when "01" & x"770" => data <= x"e5";
            when "01" & x"771" => data <= x"fe";
            when "01" & x"772" => data <= x"4c";
            when "01" & x"773" => data <= x"37";
            when "01" & x"774" => data <= x"97";
            when "01" & x"775" => data <= x"20";
            when "01" & x"776" => data <= x"28";
            when "01" & x"777" => data <= x"97";
            when "01" & x"778" => data <= x"81";
            when "01" & x"779" => data <= x"b8";
            when "01" & x"77a" => data <= x"4c";
            when "01" & x"77b" => data <= x"37";
            when "01" & x"77c" => data <= x"97";
            when "01" & x"77d" => data <= x"20";
            when "01" & x"77e" => data <= x"85";
            when "01" & x"77f" => data <= x"97";
            when "01" & x"780" => data <= x"20";
            when "01" & x"781" => data <= x"aa";
            when "01" & x"782" => data <= x"91";
            when "01" & x"783" => data <= x"18";
            when "01" & x"784" => data <= x"60";
            when "01" & x"785" => data <= x"2c";
            when "01" & x"786" => data <= x"81";
            when "01" & x"787" => data <= x"10";
            when "01" & x"788" => data <= x"10";
            when "01" & x"789" => data <= x"06";
            when "01" & x"78a" => data <= x"ad";
            when "01" & x"78b" => data <= x"e5";
            when "01" & x"78c" => data <= x"fe";
            when "01" & x"78d" => data <= x"4c";
            when "01" & x"78e" => data <= x"37";
            when "01" & x"78f" => data <= x"97";
            when "01" & x"790" => data <= x"20";
            when "01" & x"791" => data <= x"28";
            when "01" & x"792" => data <= x"97";
            when "01" & x"793" => data <= x"a1";
            when "01" & x"794" => data <= x"b8";
            when "01" & x"795" => data <= x"4c";
            when "01" & x"796" => data <= x"37";
            when "01" & x"797" => data <= x"97";
            when "01" & x"798" => data <= x"2c";
            when "01" & x"799" => data <= x"c8";
            when "01" & x"79a" => data <= x"10";
            when "01" & x"79b" => data <= x"30";
            when "01" & x"79c" => data <= x"03";
            when "01" & x"79d" => data <= x"ce";
            when "01" & x"79e" => data <= x"c8";
            when "01" & x"79f" => data <= x"10";
            when "01" & x"7a0" => data <= x"60";
            when "01" & x"7a1" => data <= x"20";
            when "01" & x"7a2" => data <= x"5a";
            when "01" & x"7a3" => data <= x"98";
            when "01" & x"7a4" => data <= x"20";
            when "01" & x"7a5" => data <= x"7e";
            when "01" & x"7a6" => data <= x"83";
            when "01" & x"7a7" => data <= x"a9";
            when "01" & x"7a8" => data <= x"01";
            when "01" & x"7a9" => data <= x"60";
            when "01" & x"7aa" => data <= x"20";
            when "01" & x"7ab" => data <= x"37";
            when "01" & x"7ac" => data <= x"98";
            when "01" & x"7ad" => data <= x"20";
            when "01" & x"7ae" => data <= x"7e";
            when "01" & x"7af" => data <= x"83";
            when "01" & x"7b0" => data <= x"20";
            when "01" & x"7b1" => data <= x"d1";
            when "01" & x"7b2" => data <= x"82";
            when "01" & x"7b3" => data <= x"90";
            when "01" & x"7b4" => data <= x"24";
            when "01" & x"7b5" => data <= x"20";
            when "01" & x"7b6" => data <= x"37";
            when "01" & x"7b7" => data <= x"98";
            when "01" & x"7b8" => data <= x"20";
            when "01" & x"7b9" => data <= x"df";
            when "01" & x"7ba" => data <= x"97";
            when "01" & x"7bb" => data <= x"20";
            when "01" & x"7bc" => data <= x"fb";
            when "01" & x"7bd" => data <= x"97";
            when "01" & x"7be" => data <= x"50";
            when "01" & x"7bf" => data <= x"16";
            when "01" & x"7c0" => data <= x"20";
            when "01" & x"7c1" => data <= x"37";
            when "01" & x"7c2" => data <= x"98";
            when "01" & x"7c3" => data <= x"20";
            when "01" & x"7c4" => data <= x"df";
            when "01" & x"7c5" => data <= x"97";
            when "01" & x"7c6" => data <= x"50";
            when "01" & x"7c7" => data <= x"11";
            when "01" & x"7c8" => data <= x"20";
            when "01" & x"7c9" => data <= x"37";
            when "01" & x"7ca" => data <= x"98";
            when "01" & x"7cb" => data <= x"20";
            when "01" & x"7cc" => data <= x"fb";
            when "01" & x"7cd" => data <= x"97";
            when "01" & x"7ce" => data <= x"50";
            when "01" & x"7cf" => data <= x"09";
            when "01" & x"7d0" => data <= x"20";
            when "01" & x"7d1" => data <= x"5a";
            when "01" & x"7d2" => data <= x"98";
            when "01" & x"7d3" => data <= x"20";
            when "01" & x"7d4" => data <= x"4f";
            when "01" & x"7d5" => data <= x"98";
            when "01" & x"7d6" => data <= x"20";
            when "01" & x"7d7" => data <= x"1e";
            when "01" & x"7d8" => data <= x"98";
            when "01" & x"7d9" => data <= x"20";
            when "01" & x"7da" => data <= x"c3";
            when "01" & x"7db" => data <= x"88";
            when "01" & x"7dc" => data <= x"a9";
            when "01" & x"7dd" => data <= x"01";
            when "01" & x"7de" => data <= x"60";
            when "01" & x"7df" => data <= x"20";
            when "01" & x"7e0" => data <= x"e1";
            when "01" & x"7e1" => data <= x"83";
            when "01" & x"7e2" => data <= x"a0";
            when "01" & x"7e3" => data <= x"02";
            when "01" & x"7e4" => data <= x"b1";
            when "01" & x"7e5" => data <= x"b0";
            when "01" & x"7e6" => data <= x"9d";
            when "01" & x"7e7" => data <= x"08";
            when "01" & x"7e8" => data <= x"0f";
            when "01" & x"7e9" => data <= x"c8";
            when "01" & x"7ea" => data <= x"b1";
            when "01" & x"7eb" => data <= x"b0";
            when "01" & x"7ec" => data <= x"9d";
            when "01" & x"7ed" => data <= x"09";
            when "01" & x"7ee" => data <= x"0f";
            when "01" & x"7ef" => data <= x"c8";
            when "01" & x"7f0" => data <= x"b1";
            when "01" & x"7f1" => data <= x"b0";
            when "01" & x"7f2" => data <= x"0a";
            when "01" & x"7f3" => data <= x"0a";
            when "01" & x"7f4" => data <= x"5d";
            when "01" & x"7f5" => data <= x"0e";
            when "01" & x"7f6" => data <= x"0f";
            when "01" & x"7f7" => data <= x"29";
            when "01" & x"7f8" => data <= x"0c";
            when "01" & x"7f9" => data <= x"10";
            when "01" & x"7fa" => data <= x"1b";
            when "01" & x"7fb" => data <= x"20";
            when "01" & x"7fc" => data <= x"e1";
            when "01" & x"7fd" => data <= x"83";
            when "01" & x"7fe" => data <= x"a0";
            when "01" & x"7ff" => data <= x"06";
            when "01" & x"800" => data <= x"b1";
            when "01" & x"801" => data <= x"b0";
            when "01" & x"802" => data <= x"9d";
            when "01" & x"803" => data <= x"0a";
            when "01" & x"804" => data <= x"0f";
            when "01" & x"805" => data <= x"c8";
            when "01" & x"806" => data <= x"b1";
            when "01" & x"807" => data <= x"b0";
            when "01" & x"808" => data <= x"9d";
            when "01" & x"809" => data <= x"0b";
            when "01" & x"80a" => data <= x"0f";
            when "01" & x"80b" => data <= x"c8";
            when "01" & x"80c" => data <= x"b1";
            when "01" & x"80d" => data <= x"b0";
            when "01" & x"80e" => data <= x"6a";
            when "01" & x"80f" => data <= x"6a";
            when "01" & x"810" => data <= x"6a";
            when "01" & x"811" => data <= x"5d";
            when "01" & x"812" => data <= x"0e";
            when "01" & x"813" => data <= x"0f";
            when "01" & x"814" => data <= x"29";
            when "01" & x"815" => data <= x"c0";
            when "01" & x"816" => data <= x"5d";
            when "01" & x"817" => data <= x"0e";
            when "01" & x"818" => data <= x"0f";
            when "01" & x"819" => data <= x"9d";
            when "01" & x"81a" => data <= x"0e";
            when "01" & x"81b" => data <= x"0f";
            when "01" & x"81c" => data <= x"b8";
            when "01" & x"81d" => data <= x"60";
            when "01" & x"81e" => data <= x"20";
            when "01" & x"81f" => data <= x"e1";
            when "01" & x"820" => data <= x"83";
            when "01" & x"821" => data <= x"a0";
            when "01" & x"822" => data <= x"0e";
            when "01" & x"823" => data <= x"b1";
            when "01" & x"824" => data <= x"b0";
            when "01" & x"825" => data <= x"29";
            when "01" & x"826" => data <= x"0a";
            when "01" & x"827" => data <= x"f0";
            when "01" & x"828" => data <= x"02";
            when "01" & x"829" => data <= x"a9";
            when "01" & x"82a" => data <= x"80";
            when "01" & x"82b" => data <= x"5d";
            when "01" & x"82c" => data <= x"0f";
            when "01" & x"82d" => data <= x"0e";
            when "01" & x"82e" => data <= x"29";
            when "01" & x"82f" => data <= x"80";
            when "01" & x"830" => data <= x"5d";
            when "01" & x"831" => data <= x"0f";
            when "01" & x"832" => data <= x"0e";
            when "01" & x"833" => data <= x"9d";
            when "01" & x"834" => data <= x"0f";
            when "01" & x"835" => data <= x"0e";
            when "01" & x"836" => data <= x"60";
            when "01" & x"837" => data <= x"20";
            when "01" & x"838" => data <= x"64";
            when "01" & x"839" => data <= x"98";
            when "01" & x"83a" => data <= x"90";
            when "01" & x"83b" => data <= x"23";
            when "01" & x"83c" => data <= x"b9";
            when "01" & x"83d" => data <= x"0f";
            when "01" & x"83e" => data <= x"0e";
            when "01" & x"83f" => data <= x"10";
            when "01" & x"840" => data <= x"22";
            when "01" & x"841" => data <= x"20";
            when "01" & x"842" => data <= x"2b";
            when "01" & x"843" => data <= x"80";
            when "01" & x"844" => data <= x"c3";
            when "01" & x"845" => data <= x"6c";
            when "01" & x"846" => data <= x"6f";
            when "01" & x"847" => data <= x"63";
            when "01" & x"848" => data <= x"6b";
            when "01" & x"849" => data <= x"65";
            when "01" & x"84a" => data <= x"64";
            when "01" & x"84b" => data <= x"00";
            when "01" & x"84c" => data <= x"20";
            when "01" & x"84d" => data <= x"3c";
            when "01" & x"84e" => data <= x"98";
            when "01" & x"84f" => data <= x"20";
            when "01" & x"850" => data <= x"e1";
            when "01" & x"851" => data <= x"83";
            when "01" & x"852" => data <= x"20";
            when "01" & x"853" => data <= x"9e";
            when "01" & x"854" => data <= x"8f";
            when "01" & x"855" => data <= x"90";
            when "01" & x"856" => data <= x"21";
            when "01" & x"857" => data <= x"4c";
            when "01" & x"858" => data <= x"02";
            when "01" & x"859" => data <= x"8f";
            when "01" & x"85a" => data <= x"20";
            when "01" & x"85b" => data <= x"64";
            when "01" & x"85c" => data <= x"98";
            when "01" & x"85d" => data <= x"b0";
            when "01" & x"85e" => data <= x"19";
            when "01" & x"85f" => data <= x"68";
            when "01" & x"860" => data <= x"68";
            when "01" & x"861" => data <= x"a9";
            when "01" & x"862" => data <= x"00";
            when "01" & x"863" => data <= x"60";
            when "01" & x"864" => data <= x"20";
            when "01" & x"865" => data <= x"06";
            when "01" & x"866" => data <= x"81";
            when "01" & x"867" => data <= x"20";
            when "01" & x"868" => data <= x"96";
            when "01" & x"869" => data <= x"82";
            when "01" & x"86a" => data <= x"90";
            when "01" & x"86b" => data <= x"0c";
            when "01" & x"86c" => data <= x"98";
            when "01" & x"86d" => data <= x"aa";
            when "01" & x"86e" => data <= x"ad";
            when "01" & x"86f" => data <= x"dc";
            when "01" & x"870" => data <= x"10";
            when "01" & x"871" => data <= x"85";
            when "01" & x"872" => data <= x"b0";
            when "01" & x"873" => data <= x"ad";
            when "01" & x"874" => data <= x"dd";
            when "01" & x"875" => data <= x"10";
            when "01" & x"876" => data <= x"85";
            when "01" & x"877" => data <= x"b1";
            when "01" & x"878" => data <= x"60";
            when "01" & x"879" => data <= x"a9";
            when "01" & x"87a" => data <= x"83";
            when "01" & x"87b" => data <= x"20";
            when "01" & x"87c" => data <= x"f4";
            when "01" & x"87d" => data <= x"ff";
            when "01" & x"87e" => data <= x"8c";
            when "01" & x"87f" => data <= x"d0";
            when "01" & x"880" => data <= x"10";
            when "01" & x"881" => data <= x"a9";
            when "01" & x"882" => data <= x"84";
            when "01" & x"883" => data <= x"20";
            when "01" & x"884" => data <= x"f4";
            when "01" & x"885" => data <= x"ff";
            when "01" & x"886" => data <= x"98";
            when "01" & x"887" => data <= x"38";
            when "01" & x"888" => data <= x"ed";
            when "01" & x"889" => data <= x"d0";
            when "01" & x"88a" => data <= x"10";
            when "01" & x"88b" => data <= x"8d";
            when "01" & x"88c" => data <= x"d1";
            when "01" & x"88d" => data <= x"10";
            when "01" & x"88e" => data <= x"60";
            when "01" & x"88f" => data <= x"a2";
            when "01" & x"890" => data <= x"0a";
            when "01" & x"891" => data <= x"20";
            when "01" & x"892" => data <= x"2c";
            when "01" & x"893" => data <= x"99";
            when "01" & x"894" => data <= x"20";
            when "01" & x"895" => data <= x"9e";
            when "01" & x"896" => data <= x"98";
            when "01" & x"897" => data <= x"a0";
            when "01" & x"898" => data <= x"d5";
            when "01" & x"899" => data <= x"a9";
            when "01" & x"89a" => data <= x"ff";
            when "01" & x"89b" => data <= x"91";
            when "01" & x"89c" => data <= x"b0";
            when "01" & x"89d" => data <= x"60";
            when "01" & x"89e" => data <= x"48";
            when "01" & x"89f" => data <= x"a6";
            when "01" & x"8a0" => data <= x"f4";
            when "01" & x"8a1" => data <= x"a9";
            when "01" & x"8a2" => data <= x"00";
            when "01" & x"8a3" => data <= x"85";
            when "01" & x"8a4" => data <= x"b0";
            when "01" & x"8a5" => data <= x"bd";
            when "01" & x"8a6" => data <= x"f0";
            when "01" & x"8a7" => data <= x"0d";
            when "01" & x"8a8" => data <= x"85";
            when "01" & x"8a9" => data <= x"b1";
            when "01" & x"8aa" => data <= x"68";
            when "01" & x"8ab" => data <= x"60";
            when "01" & x"8ac" => data <= x"00";
            when "01" & x"8ad" => data <= x"00";
            when "01" & x"8ae" => data <= x"00";
            when "01" & x"8af" => data <= x"00";
            when "01" & x"8b0" => data <= x"00";
            when "01" & x"8b1" => data <= x"00";
            when "01" & x"8b2" => data <= x"00";
            when "01" & x"8b3" => data <= x"00";
            when "01" & x"8b4" => data <= x"00";
            when "01" & x"8b5" => data <= x"00";
            when "01" & x"8b6" => data <= x"00";
            when "01" & x"8b7" => data <= x"00";
            when "01" & x"8b8" => data <= x"00";
            when "01" & x"8b9" => data <= x"00";
            when "01" & x"8ba" => data <= x"00";
            when "01" & x"8bb" => data <= x"00";
            when "01" & x"8bc" => data <= x"00";
            when "01" & x"8bd" => data <= x"00";
            when "01" & x"8be" => data <= x"00";
            when "01" & x"8bf" => data <= x"00";
            when "01" & x"8c0" => data <= x"00";
            when "01" & x"8c1" => data <= x"00";
            when "01" & x"8c2" => data <= x"00";
            when "01" & x"8c3" => data <= x"00";
            when "01" & x"8c4" => data <= x"00";
            when "01" & x"8c5" => data <= x"00";
            when "01" & x"8c6" => data <= x"00";
            when "01" & x"8c7" => data <= x"00";
            when "01" & x"8c8" => data <= x"00";
            when "01" & x"8c9" => data <= x"00";
            when "01" & x"8ca" => data <= x"00";
            when "01" & x"8cb" => data <= x"00";
            when "01" & x"8cc" => data <= x"00";
            when "01" & x"8cd" => data <= x"00";
            when "01" & x"8ce" => data <= x"00";
            when "01" & x"8cf" => data <= x"00";
            when "01" & x"8d0" => data <= x"00";
            when "01" & x"8d1" => data <= x"00";
            when "01" & x"8d2" => data <= x"00";
            when "01" & x"8d3" => data <= x"00";
            when "01" & x"8d4" => data <= x"00";
            when "01" & x"8d5" => data <= x"00";
            when "01" & x"8d6" => data <= x"00";
            when "01" & x"8d7" => data <= x"00";
            when "01" & x"8d8" => data <= x"00";
            when "01" & x"8d9" => data <= x"00";
            when "01" & x"8da" => data <= x"00";
            when "01" & x"8db" => data <= x"00";
            when "01" & x"8dc" => data <= x"00";
            when "01" & x"8dd" => data <= x"00";
            when "01" & x"8de" => data <= x"00";
            when "01" & x"8df" => data <= x"00";
            when "01" & x"8e0" => data <= x"00";
            when "01" & x"8e1" => data <= x"00";
            when "01" & x"8e2" => data <= x"00";
            when "01" & x"8e3" => data <= x"00";
            when "01" & x"8e4" => data <= x"00";
            when "01" & x"8e5" => data <= x"00";
            when "01" & x"8e6" => data <= x"00";
            when "01" & x"8e7" => data <= x"00";
            when "01" & x"8e8" => data <= x"00";
            when "01" & x"8e9" => data <= x"00";
            when "01" & x"8ea" => data <= x"00";
            when "01" & x"8eb" => data <= x"00";
            when "01" & x"8ec" => data <= x"00";
            when "01" & x"8ed" => data <= x"00";
            when "01" & x"8ee" => data <= x"00";
            when "01" & x"8ef" => data <= x"00";
            when "01" & x"8f0" => data <= x"00";
            when "01" & x"8f1" => data <= x"00";
            when "01" & x"8f2" => data <= x"00";
            when "01" & x"8f3" => data <= x"00";
            when "01" & x"8f4" => data <= x"00";
            when "01" & x"8f5" => data <= x"00";
            when "01" & x"8f6" => data <= x"00";
            when "01" & x"8f7" => data <= x"00";
            when "01" & x"8f8" => data <= x"00";
            when "01" & x"8f9" => data <= x"00";
            when "01" & x"8fa" => data <= x"00";
            when "01" & x"8fb" => data <= x"00";
            when "01" & x"8fc" => data <= x"00";
            when "01" & x"8fd" => data <= x"00";
            when "01" & x"8fe" => data <= x"00";
            when "01" & x"8ff" => data <= x"00";
            when "01" & x"900" => data <= x"00";
            when "01" & x"901" => data <= x"00";
            when "01" & x"902" => data <= x"00";
            when "01" & x"903" => data <= x"00";
            when "01" & x"904" => data <= x"00";
            when "01" & x"905" => data <= x"60";
            when "01" & x"906" => data <= x"20";
            when "01" & x"907" => data <= x"e1";
            when "01" & x"908" => data <= x"83";
            when "01" & x"909" => data <= x"a9";
            when "01" & x"90a" => data <= x"0f";
            when "01" & x"90b" => data <= x"a2";
            when "01" & x"90c" => data <= x"01";
            when "01" & x"90d" => data <= x"a0";
            when "01" & x"90e" => data <= x"00";
            when "01" & x"90f" => data <= x"f0";
            when "01" & x"910" => data <= x"25";
            when "01" & x"911" => data <= x"a9";
            when "01" & x"912" => data <= x"c7";
            when "01" & x"913" => data <= x"a2";
            when "01" & x"914" => data <= x"00";
            when "01" & x"915" => data <= x"f0";
            when "01" & x"916" => data <= x"f6";
            when "01" & x"917" => data <= x"aa";
            when "01" & x"918" => data <= x"a9";
            when "01" & x"919" => data <= x"03";
            when "01" & x"91a" => data <= x"d0";
            when "01" & x"91b" => data <= x"1a";
            when "01" & x"91c" => data <= x"a9";
            when "01" & x"91d" => data <= x"ec";
            when "01" & x"91e" => data <= x"d0";
            when "01" & x"91f" => data <= x"12";
            when "01" & x"920" => data <= x"a9";
            when "01" & x"921" => data <= x"c7";
            when "01" & x"922" => data <= x"d0";
            when "01" & x"923" => data <= x"0e";
            when "01" & x"924" => data <= x"a9";
            when "01" & x"925" => data <= x"ea";
            when "01" & x"926" => data <= x"d0";
            when "01" & x"927" => data <= x"0a";
            when "01" & x"928" => data <= x"a9";
            when "01" & x"929" => data <= x"a8";
            when "01" & x"92a" => data <= x"d0";
            when "01" & x"92b" => data <= x"06";
            when "01" & x"92c" => data <= x"a9";
            when "01" & x"92d" => data <= x"8f";
            when "01" & x"92e" => data <= x"d0";
            when "01" & x"92f" => data <= x"06";
            when "01" & x"930" => data <= x"a9";
            when "01" & x"931" => data <= x"ff";
            when "01" & x"932" => data <= x"a2";
            when "01" & x"933" => data <= x"00";
            when "01" & x"934" => data <= x"a0";
            when "01" & x"935" => data <= x"ff";
            when "01" & x"936" => data <= x"4c";
            when "01" & x"937" => data <= x"f4";
            when "01" & x"938" => data <= x"ff";
            when "01" & x"939" => data <= x"4c";
            when "01" & x"93a" => data <= x"2e";
            when "01" & x"93b" => data <= x"21";
            when "01" & x"93c" => data <= x"42";
            when "01" & x"93d" => data <= x"4f";
            when "01" & x"93e" => data <= x"4f";
            when "01" & x"93f" => data <= x"54";
            when "01" & x"940" => data <= x"0d";
            when "01" & x"941" => data <= x"45";
            when "01" & x"942" => data <= x"2e";
            when "01" & x"943" => data <= x"21";
            when "01" & x"944" => data <= x"42";
            when "01" & x"945" => data <= x"4f";
            when "01" & x"946" => data <= x"4f";
            when "01" & x"947" => data <= x"54";
            when "01" & x"948" => data <= x"0d";
            when "01" & x"949" => data <= x"1b";
            when "01" & x"94a" => data <= x"ff";
            when "01" & x"94b" => data <= x"1e";
            when "01" & x"94c" => data <= x"ff";
            when "01" & x"94d" => data <= x"21";
            when "01" & x"94e" => data <= x"ff";
            when "01" & x"94f" => data <= x"24";
            when "01" & x"950" => data <= x"ff";
            when "01" & x"951" => data <= x"27";
            when "01" & x"952" => data <= x"ff";
            when "01" & x"953" => data <= x"2a";
            when "01" & x"954" => data <= x"ff";
            when "01" & x"955" => data <= x"2d";
            when "01" & x"956" => data <= x"ff";
            when "01" & x"957" => data <= x"7b";
            when "01" & x"958" => data <= x"95";
            when "01" & x"959" => data <= x"00";
            when "01" & x"95a" => data <= x"07";
            when "01" & x"95b" => data <= x"90";
            when "01" & x"95c" => data <= x"00";
            when "01" & x"95d" => data <= x"c1";
            when "01" & x"95e" => data <= x"90";
            when "01" & x"95f" => data <= x"00";
            when "01" & x"960" => data <= x"aa";
            when "01" & x"961" => data <= x"91";
            when "01" & x"962" => data <= x"00";
            when "01" & x"963" => data <= x"d0";
            when "01" & x"964" => data <= x"95";
            when "01" & x"965" => data <= x"00";
            when "01" & x"966" => data <= x"93";
            when "01" & x"967" => data <= x"8e";
            when "01" & x"968" => data <= x"00";
            when "01" & x"969" => data <= x"aa";
            when "01" & x"96a" => data <= x"95";
            when "01" & x"96b" => data <= x"00";
            when "01" & x"96c" => data <= x"1b";
            when "01" & x"96d" => data <= x"8c";
            when "01" & x"96e" => data <= x"d3";
            when "01" & x"96f" => data <= x"6b";
            when "01" & x"970" => data <= x"d3";
            when "01" & x"971" => data <= x"1d";
            when "01" & x"972" => data <= x"e1";
            when "01" & x"973" => data <= x"dc";
            when "01" & x"974" => data <= x"97";
            when "01" & x"975" => data <= x"89";
            when "01" & x"976" => data <= x"90";
            when "01" & x"977" => data <= x"87";
            when "01" & x"978" => data <= x"86";
            when "01" & x"979" => data <= x"87";
            when "01" & x"97a" => data <= x"84";
            when "01" & x"97b" => data <= x"8d";
            when "01" & x"97c" => data <= x"8d";
            when "01" & x"97d" => data <= x"97";
            when "01" & x"97e" => data <= x"f1";
            when "01" & x"97f" => data <= x"3c";
            when "01" & x"980" => data <= x"bc";
            when "01" & x"981" => data <= x"8f";
            when "01" & x"982" => data <= x"9b";
            when "01" & x"983" => data <= x"95";
            when "01" & x"984" => data <= x"93";
            when "01" & x"985" => data <= x"85";
            when "01" & x"986" => data <= x"b4";
            when "01" & x"987" => data <= x"bf";
            when "01" & x"988" => data <= x"c7";
            when "01" & x"989" => data <= x"cf";
            when "01" & x"98a" => data <= x"a0";
            when "01" & x"98b" => data <= x"a9";
            when "01" & x"98c" => data <= x"87";
            when "01" & x"98d" => data <= x"87";
            when "01" & x"98e" => data <= x"97";
            when "01" & x"98f" => data <= x"97";
            when "01" & x"990" => data <= x"97";
            when "01" & x"991" => data <= x"97";
            when "01" & x"992" => data <= x"97";
            when "01" & x"993" => data <= x"97";
            when "01" & x"994" => data <= x"12";
            when "01" & x"995" => data <= x"32";
            when "01" & x"996" => data <= x"5d";
            when "01" & x"997" => data <= x"cd";
            when "01" & x"998" => data <= x"a2";
            when "01" & x"999" => data <= x"bd";
            when "01" & x"99a" => data <= x"87";
            when "01" & x"99b" => data <= x"8d";
            when "01" & x"99c" => data <= x"8d";
            when "01" & x"99d" => data <= x"8d";
            when "01" & x"99e" => data <= x"8d";
            when "01" & x"99f" => data <= x"8d";
            when "01" & x"9a0" => data <= x"8d";
            when "01" & x"9a1" => data <= x"8d";
            when "01" & x"9a2" => data <= x"74";
            when "01" & x"9a3" => data <= x"54";
            when "01" & x"9a4" => data <= x"00";
            when "01" & x"9a5" => data <= x"0f";
            when "01" & x"9a6" => data <= x"1a";
            when "01" & x"9a7" => data <= x"0f";
            when "01" & x"9a8" => data <= x"1a";
            when "01" & x"9a9" => data <= x"63";
            when "01" & x"9aa" => data <= x"43";
            when "01" & x"9ab" => data <= x"b7";
            when "01" & x"9ac" => data <= x"7d";
            when "01" & x"9ad" => data <= x"7d";
            when "01" & x"9ae" => data <= x"65";
            when "01" & x"9af" => data <= x"65";
            when "01" & x"9b0" => data <= x"cf";
            when "01" & x"9b1" => data <= x"00";
            when "01" & x"9b2" => data <= x"14";
            when "01" & x"9b3" => data <= x"83";
            when "01" & x"9b4" => data <= x"85";
            when "01" & x"9b5" => data <= x"97";
            when "01" & x"9b6" => data <= x"97";
            when "01" & x"9b7" => data <= x"97";
            when "01" & x"9b8" => data <= x"97";
            when "01" & x"9b9" => data <= x"96";
            when "01" & x"9ba" => data <= x"97";
            when "01" & x"9bb" => data <= x"97";
            when "01" & x"9bc" => data <= x"96";
            when "01" & x"9bd" => data <= x"04";
            when "01" & x"9be" => data <= x"02";
            when "01" & x"9bf" => data <= x"03";
            when "01" & x"9c0" => data <= x"06";
            when "01" & x"9c1" => data <= x"07";
            when "01" & x"9c2" => data <= x"04";
            when "01" & x"9c3" => data <= x"04";
            when "01" & x"9c4" => data <= x"04";
            when "01" & x"9c5" => data <= x"04";
            when "01" & x"9c6" => data <= x"98";
            when "01" & x"9c7" => data <= x"a2";
            when "01" & x"9c8" => data <= x"ff";
            when "01" & x"9c9" => data <= x"a0";
            when "01" & x"9ca" => data <= x"0e";
            when "01" & x"9cb" => data <= x"48";
            when "01" & x"9cc" => data <= x"20";
            when "01" & x"9cd" => data <= x"65";
            when "01" & x"9ce" => data <= x"80";
            when "01" & x"9cf" => data <= x"0d";
            when "01" & x"9d0" => data <= x"44";
            when "01" & x"9d1" => data <= x"46";
            when "01" & x"9d2" => data <= x"53";
            when "01" & x"9d3" => data <= x"20";
            when "01" & x"9d4" => data <= x"30";
            when "01" & x"9d5" => data <= x"2e";
            when "01" & x"9d6" => data <= x"39";
            when "01" & x"9d7" => data <= x"30";
            when "01" & x"9d8" => data <= x"0d";
            when "01" & x"9d9" => data <= x"86";
            when "01" & x"9da" => data <= x"b8";
            when "01" & x"9db" => data <= x"20";
            when "01" & x"9dc" => data <= x"cb";
            when "01" & x"9dd" => data <= x"9f";
            when "01" & x"9de" => data <= x"20";
            when "01" & x"9df" => data <= x"19";
            when "01" & x"9e0" => data <= x"9a";
            when "01" & x"9e1" => data <= x"20";
            when "01" & x"9e2" => data <= x"9a";
            when "01" & x"9e3" => data <= x"9f";
            when "01" & x"9e4" => data <= x"88";
            when "01" & x"9e5" => data <= x"d0";
            when "01" & x"9e6" => data <= x"f4";
            when "01" & x"9e7" => data <= x"68";
            when "01" & x"9e8" => data <= x"a8";
            when "01" & x"9e9" => data <= x"a2";
            when "01" & x"9ea" => data <= x"a0";
            when "01" & x"9eb" => data <= x"4c";
            when "01" & x"9ec" => data <= x"71";
            when "01" & x"9ed" => data <= x"86";
            when "01" & x"9ee" => data <= x"98";
            when "01" & x"9ef" => data <= x"a2";
            when "01" & x"9f0" => data <= x"74";
            when "01" & x"9f1" => data <= x"a0";
            when "01" & x"9f2" => data <= x"05";
            when "01" & x"9f3" => data <= x"d0";
            when "01" & x"9f4" => data <= x"d6";
            when "01" & x"9f5" => data <= x"20";
            when "01" & x"9f6" => data <= x"bf";
            when "01" & x"9f7" => data <= x"86";
            when "01" & x"9f8" => data <= x"f0";
            when "01" & x"9f9" => data <= x"60";
            when "01" & x"9fa" => data <= x"20";
            when "01" & x"9fb" => data <= x"c5";
            when "01" & x"9fc" => data <= x"ff";
            when "01" & x"9fd" => data <= x"90";
            when "01" & x"9fe" => data <= x"fb";
            when "01" & x"9ff" => data <= x"b0";
            when "01" & x"a00" => data <= x"e8";
            when "01" & x"a01" => data <= x"20";
            when "01" & x"a02" => data <= x"bf";
            when "01" & x"a03" => data <= x"86";
            when "01" & x"a04" => data <= x"d0";
            when "01" & x"a05" => data <= x"54";
            when "01" & x"a06" => data <= x"20";
            when "01" & x"a07" => data <= x"33";
            when "01" & x"a08" => data <= x"80";
            when "01" & x"a09" => data <= x"dc";
            when "01" & x"a0a" => data <= x"53";
            when "01" & x"a0b" => data <= x"79";
            when "01" & x"a0c" => data <= x"6e";
            when "01" & x"a0d" => data <= x"74";
            when "01" & x"a0e" => data <= x"61";
            when "01" & x"a0f" => data <= x"78";
            when "01" & x"a10" => data <= x"3a";
            when "01" & x"a11" => data <= x"20";
            when "01" & x"a12" => data <= x"ea";
            when "01" & x"a13" => data <= x"20";
            when "01" & x"a14" => data <= x"19";
            when "01" & x"a15" => data <= x"9a";
            when "01" & x"a16" => data <= x"4c";
            when "01" & x"a17" => data <= x"8a";
            when "01" & x"a18" => data <= x"80";
            when "01" & x"a19" => data <= x"a6";
            when "01" & x"a1a" => data <= x"b8";
            when "01" & x"a1b" => data <= x"e8";
            when "01" & x"a1c" => data <= x"bd";
            when "01" & x"a1d" => data <= x"b8";
            when "01" & x"a1e" => data <= x"85";
            when "01" & x"a1f" => data <= x"30";
            when "01" & x"a20" => data <= x"06";
            when "01" & x"a21" => data <= x"20";
            when "01" & x"a22" => data <= x"9c";
            when "01" & x"a23" => data <= x"80";
            when "01" & x"a24" => data <= x"4c";
            when "01" & x"a25" => data <= x"1b";
            when "01" & x"a26" => data <= x"9a";
            when "01" & x"a27" => data <= x"e8";
            when "01" & x"a28" => data <= x"e8";
            when "01" & x"a29" => data <= x"86";
            when "01" & x"a2a" => data <= x"b8";
            when "01" & x"a2b" => data <= x"bd";
            when "01" & x"a2c" => data <= x"b8";
            when "01" & x"a2d" => data <= x"85";
            when "01" & x"a2e" => data <= x"20";
            when "01" & x"a2f" => data <= x"34";
            when "01" & x"a30" => data <= x"9a";
            when "01" & x"a31" => data <= x"20";
            when "01" & x"a32" => data <= x"05";
            when "01" & x"a33" => data <= x"82";
            when "01" & x"a34" => data <= x"20";
            when "01" & x"a35" => data <= x"e1";
            when "01" & x"a36" => data <= x"83";
            when "01" & x"a37" => data <= x"29";
            when "01" & x"a38" => data <= x"0f";
            when "01" & x"a39" => data <= x"f0";
            when "01" & x"a3a" => data <= x"1f";
            when "01" & x"a3b" => data <= x"a8";
            when "01" & x"a3c" => data <= x"a9";
            when "01" & x"a3d" => data <= x"20";
            when "01" & x"a3e" => data <= x"20";
            when "01" & x"a3f" => data <= x"9c";
            when "01" & x"a40" => data <= x"80";
            when "01" & x"a41" => data <= x"a2";
            when "01" & x"a42" => data <= x"00";
            when "01" & x"a43" => data <= x"bd";
            when "01" & x"a44" => data <= x"5b";
            when "01" & x"a45" => data <= x"9a";
            when "01" & x"a46" => data <= x"f0";
            when "01" & x"a47" => data <= x"03";
            when "01" & x"a48" => data <= x"e8";
            when "01" & x"a49" => data <= x"d0";
            when "01" & x"a4a" => data <= x"f8";
            when "01" & x"a4b" => data <= x"88";
            when "01" & x"a4c" => data <= x"d0";
            when "01" & x"a4d" => data <= x"fa";
            when "01" & x"a4e" => data <= x"e8";
            when "01" & x"a4f" => data <= x"bd";
            when "01" & x"a50" => data <= x"5b";
            when "01" & x"a51" => data <= x"9a";
            when "01" & x"a52" => data <= x"f0";
            when "01" & x"a53" => data <= x"06";
            when "01" & x"a54" => data <= x"20";
            when "01" & x"a55" => data <= x"9c";
            when "01" & x"a56" => data <= x"80";
            when "01" & x"a57" => data <= x"4c";
            when "01" & x"a58" => data <= x"4e";
            when "01" & x"a59" => data <= x"9a";
            when "01" & x"a5a" => data <= x"60";
            when "01" & x"a5b" => data <= x"00";
            when "01" & x"a5c" => data <= x"3c";
            when "01" & x"a5d" => data <= x"66";
            when "01" & x"a5e" => data <= x"73";
            when "01" & x"a5f" => data <= x"70";
            when "01" & x"a60" => data <= x"3e";
            when "01" & x"a61" => data <= x"00";
            when "01" & x"a62" => data <= x"3c";
            when "01" & x"a63" => data <= x"61";
            when "01" & x"a64" => data <= x"66";
            when "01" & x"a65" => data <= x"73";
            when "01" & x"a66" => data <= x"70";
            when "01" & x"a67" => data <= x"3e";
            when "01" & x"a68" => data <= x"00";
            when "01" & x"a69" => data <= x"28";
            when "01" & x"a6a" => data <= x"4c";
            when "01" & x"a6b" => data <= x"29";
            when "01" & x"a6c" => data <= x"00";
            when "01" & x"a6d" => data <= x"3c";
            when "01" & x"a6e" => data <= x"73";
            when "01" & x"a6f" => data <= x"72";
            when "01" & x"a70" => data <= x"63";
            when "01" & x"a71" => data <= x"20";
            when "01" & x"a72" => data <= x"64";
            when "01" & x"a73" => data <= x"72";
            when "01" & x"a74" => data <= x"76";
            when "01" & x"a75" => data <= x"3e";
            when "01" & x"a76" => data <= x"00";
            when "01" & x"a77" => data <= x"3c";
            when "01" & x"a78" => data <= x"64";
            when "01" & x"a79" => data <= x"65";
            when "01" & x"a7a" => data <= x"73";
            when "01" & x"a7b" => data <= x"74";
            when "01" & x"a7c" => data <= x"20";
            when "01" & x"a7d" => data <= x"64";
            when "01" & x"a7e" => data <= x"72";
            when "01" & x"a7f" => data <= x"76";
            when "01" & x"a80" => data <= x"3e";
            when "01" & x"a81" => data <= x"00";
            when "01" & x"a82" => data <= x"3c";
            when "01" & x"a83" => data <= x"64";
            when "01" & x"a84" => data <= x"65";
            when "01" & x"a85" => data <= x"73";
            when "01" & x"a86" => data <= x"74";
            when "01" & x"a87" => data <= x"20";
            when "01" & x"a88" => data <= x"64";
            when "01" & x"a89" => data <= x"72";
            when "01" & x"a8a" => data <= x"76";
            when "01" & x"a8b" => data <= x"3e";
            when "01" & x"a8c" => data <= x"20";
            when "01" & x"a8d" => data <= x"3c";
            when "01" & x"a8e" => data <= x"61";
            when "01" & x"a8f" => data <= x"66";
            when "01" & x"a90" => data <= x"73";
            when "01" & x"a91" => data <= x"70";
            when "01" & x"a92" => data <= x"3e";
            when "01" & x"a93" => data <= x"00";
            when "01" & x"a94" => data <= x"3c";
            when "01" & x"a95" => data <= x"6f";
            when "01" & x"a96" => data <= x"6c";
            when "01" & x"a97" => data <= x"64";
            when "01" & x"a98" => data <= x"20";
            when "01" & x"a99" => data <= x"66";
            when "01" & x"a9a" => data <= x"73";
            when "01" & x"a9b" => data <= x"70";
            when "01" & x"a9c" => data <= x"3e";
            when "01" & x"a9d" => data <= x"00";
            when "01" & x"a9e" => data <= x"3c";
            when "01" & x"a9f" => data <= x"6e";
            when "01" & x"aa0" => data <= x"65";
            when "01" & x"aa1" => data <= x"77";
            when "01" & x"aa2" => data <= x"20";
            when "01" & x"aa3" => data <= x"66";
            when "01" & x"aa4" => data <= x"73";
            when "01" & x"aa5" => data <= x"70";
            when "01" & x"aa6" => data <= x"3e";
            when "01" & x"aa7" => data <= x"00";
            when "01" & x"aa8" => data <= x"28";
            when "01" & x"aa9" => data <= x"3c";
            when "01" & x"aaa" => data <= x"64";
            when "01" & x"aab" => data <= x"69";
            when "01" & x"aac" => data <= x"72";
            when "01" & x"aad" => data <= x"3e";
            when "01" & x"aae" => data <= x"29";
            when "01" & x"aaf" => data <= x"00";
            when "01" & x"ab0" => data <= x"28";
            when "01" & x"ab1" => data <= x"3c";
            when "01" & x"ab2" => data <= x"64";
            when "01" & x"ab3" => data <= x"72";
            when "01" & x"ab4" => data <= x"76";
            when "01" & x"ab5" => data <= x"3e";
            when "01" & x"ab6" => data <= x"29";
            when "01" & x"ab7" => data <= x"00";
            when "01" & x"ab8" => data <= x"3c";
            when "01" & x"ab9" => data <= x"74";
            when "01" & x"aba" => data <= x"69";
            when "01" & x"abb" => data <= x"74";
            when "01" & x"abc" => data <= x"6c";
            when "01" & x"abd" => data <= x"65";
            when "01" & x"abe" => data <= x"3e";
            when "01" & x"abf" => data <= x"00";
            when "01" & x"ac0" => data <= x"20";
            when "01" & x"ac1" => data <= x"58";
            when "01" & x"ac2" => data <= x"83";
            when "01" & x"ac3" => data <= x"20";
            when "01" & x"ac4" => data <= x"65";
            when "01" & x"ac5" => data <= x"80";
            when "01" & x"ac6" => data <= x"43";
            when "01" & x"ac7" => data <= x"6f";
            when "01" & x"ac8" => data <= x"6d";
            when "01" & x"ac9" => data <= x"70";
            when "01" & x"aca" => data <= x"61";
            when "01" & x"acb" => data <= x"63";
            when "01" & x"acc" => data <= x"74";
            when "01" & x"acd" => data <= x"69";
            when "01" & x"ace" => data <= x"6e";
            when "01" & x"acf" => data <= x"67";
            when "01" & x"ad0" => data <= x"20";
            when "01" & x"ad1" => data <= x"64";
            when "01" & x"ad2" => data <= x"72";
            when "01" & x"ad3" => data <= x"69";
            when "01" & x"ad4" => data <= x"76";
            when "01" & x"ad5" => data <= x"65";
            when "01" & x"ad6" => data <= x"20";
            when "01" & x"ad7" => data <= x"8d";
            when "01" & x"ad8" => data <= x"d2";
            when "01" & x"ad9" => data <= x"10";
            when "01" & x"ada" => data <= x"8d";
            when "01" & x"adb" => data <= x"d3";
            when "01" & x"adc" => data <= x"10";
            when "01" & x"add" => data <= x"20";
            when "01" & x"ade" => data <= x"ca";
            when "01" & x"adf" => data <= x"80";
            when "01" & x"ae0" => data <= x"20";
            when "01" & x"ae1" => data <= x"9a";
            when "01" & x"ae2" => data <= x"9f";
            when "01" & x"ae3" => data <= x"a0";
            when "01" & x"ae4" => data <= x"00";
            when "01" & x"ae5" => data <= x"20";
            when "01" & x"ae6" => data <= x"05";
            when "01" & x"ae7" => data <= x"8e";
            when "01" & x"ae8" => data <= x"20";
            when "01" & x"ae9" => data <= x"79";
            when "01" & x"aea" => data <= x"98";
            when "01" & x"aeb" => data <= x"20";
            when "01" & x"aec" => data <= x"47";
            when "01" & x"aed" => data <= x"83";
            when "01" & x"aee" => data <= x"ac";
            when "01" & x"aef" => data <= x"05";
            when "01" & x"af0" => data <= x"0f";
            when "01" & x"af1" => data <= x"84";
            when "01" & x"af2" => data <= x"cc";
            when "01" & x"af3" => data <= x"a9";
            when "01" & x"af4" => data <= x"02";
            when "01" & x"af5" => data <= x"85";
            when "01" & x"af6" => data <= x"ca";
            when "01" & x"af7" => data <= x"a9";
            when "01" & x"af8" => data <= x"00";
            when "01" & x"af9" => data <= x"85";
            when "01" & x"afa" => data <= x"cb";
            when "01" & x"afb" => data <= x"a4";
            when "01" & x"afc" => data <= x"cc";
            when "01" & x"afd" => data <= x"20";
            when "01" & x"afe" => data <= x"19";
            when "01" & x"aff" => data <= x"82";
            when "01" & x"b00" => data <= x"c0";
            when "01" & x"b01" => data <= x"f8";
            when "01" & x"b02" => data <= x"d0";
            when "01" & x"b03" => data <= x"3c";
            when "01" & x"b04" => data <= x"20";
            when "01" & x"b05" => data <= x"65";
            when "01" & x"b06" => data <= x"80";
            when "01" & x"b07" => data <= x"44";
            when "01" & x"b08" => data <= x"69";
            when "01" & x"b09" => data <= x"73";
            when "01" & x"b0a" => data <= x"6b";
            when "01" & x"b0b" => data <= x"20";
            when "01" & x"b0c" => data <= x"63";
            when "01" & x"b0d" => data <= x"6f";
            when "01" & x"b0e" => data <= x"6d";
            when "01" & x"b0f" => data <= x"70";
            when "01" & x"b10" => data <= x"61";
            when "01" & x"b11" => data <= x"63";
            when "01" & x"b12" => data <= x"74";
            when "01" & x"b13" => data <= x"65";
            when "01" & x"b14" => data <= x"64";
            when "01" & x"b15" => data <= x"20";
            when "01" & x"b16" => data <= x"ea";
            when "01" & x"b17" => data <= x"38";
            when "01" & x"b18" => data <= x"ad";
            when "01" & x"b19" => data <= x"07";
            when "01" & x"b1a" => data <= x"0f";
            when "01" & x"b1b" => data <= x"e5";
            when "01" & x"b1c" => data <= x"ca";
            when "01" & x"b1d" => data <= x"48";
            when "01" & x"b1e" => data <= x"ad";
            when "01" & x"b1f" => data <= x"06";
            when "01" & x"b20" => data <= x"0f";
            when "01" & x"b21" => data <= x"29";
            when "01" & x"b22" => data <= x"03";
            when "01" & x"b23" => data <= x"e5";
            when "01" & x"b24" => data <= x"cb";
            when "01" & x"b25" => data <= x"20";
            when "01" & x"b26" => data <= x"ca";
            when "01" & x"b27" => data <= x"80";
            when "01" & x"b28" => data <= x"68";
            when "01" & x"b29" => data <= x"20";
            when "01" & x"b2a" => data <= x"c2";
            when "01" & x"b2b" => data <= x"80";
            when "01" & x"b2c" => data <= x"20";
            when "01" & x"b2d" => data <= x"65";
            when "01" & x"b2e" => data <= x"80";
            when "01" & x"b2f" => data <= x"20";
            when "01" & x"b30" => data <= x"66";
            when "01" & x"b31" => data <= x"72";
            when "01" & x"b32" => data <= x"65";
            when "01" & x"b33" => data <= x"65";
            when "01" & x"b34" => data <= x"20";
            when "01" & x"b35" => data <= x"73";
            when "01" & x"b36" => data <= x"65";
            when "01" & x"b37" => data <= x"63";
            when "01" & x"b38" => data <= x"74";
            when "01" & x"b39" => data <= x"6f";
            when "01" & x"b3a" => data <= x"72";
            when "01" & x"b3b" => data <= x"73";
            when "01" & x"b3c" => data <= x"0d";
            when "01" & x"b3d" => data <= x"a9";
            when "01" & x"b3e" => data <= x"04";
            when "01" & x"b3f" => data <= x"60";
            when "01" & x"b40" => data <= x"84";
            when "01" & x"b41" => data <= x"cc";
            when "01" & x"b42" => data <= x"20";
            when "01" & x"b43" => data <= x"fc";
            when "01" & x"b44" => data <= x"82";
            when "01" & x"b45" => data <= x"a4";
            when "01" & x"b46" => data <= x"cc";
            when "01" & x"b47" => data <= x"b9";
            when "01" & x"b48" => data <= x"0e";
            when "01" & x"b49" => data <= x"0f";
            when "01" & x"b4a" => data <= x"29";
            when "01" & x"b4b" => data <= x"30";
            when "01" & x"b4c" => data <= x"19";
            when "01" & x"b4d" => data <= x"0d";
            when "01" & x"b4e" => data <= x"0f";
            when "01" & x"b4f" => data <= x"19";
            when "01" & x"b50" => data <= x"0c";
            when "01" & x"b51" => data <= x"0f";
            when "01" & x"b52" => data <= x"f0";
            when "01" & x"b53" => data <= x"61";
            when "01" & x"b54" => data <= x"a9";
            when "01" & x"b55" => data <= x"00";
            when "01" & x"b56" => data <= x"85";
            when "01" & x"b57" => data <= x"be";
            when "01" & x"b58" => data <= x"85";
            when "01" & x"b59" => data <= x"c2";
            when "01" & x"b5a" => data <= x"a9";
            when "01" & x"b5b" => data <= x"ff";
            when "01" & x"b5c" => data <= x"18";
            when "01" & x"b5d" => data <= x"79";
            when "01" & x"b5e" => data <= x"0c";
            when "01" & x"b5f" => data <= x"0f";
            when "01" & x"b60" => data <= x"a9";
            when "01" & x"b61" => data <= x"00";
            when "01" & x"b62" => data <= x"79";
            when "01" & x"b63" => data <= x"0d";
            when "01" & x"b64" => data <= x"0f";
            when "01" & x"b65" => data <= x"85";
            when "01" & x"b66" => data <= x"c6";
            when "01" & x"b67" => data <= x"b9";
            when "01" & x"b68" => data <= x"0e";
            when "01" & x"b69" => data <= x"0f";
            when "01" & x"b6a" => data <= x"08";
            when "01" & x"b6b" => data <= x"20";
            when "01" & x"b6c" => data <= x"fd";
            when "01" & x"b6d" => data <= x"81";
            when "01" & x"b6e" => data <= x"28";
            when "01" & x"b6f" => data <= x"69";
            when "01" & x"b70" => data <= x"00";
            when "01" & x"b71" => data <= x"85";
            when "01" & x"b72" => data <= x"c7";
            when "01" & x"b73" => data <= x"b9";
            when "01" & x"b74" => data <= x"0f";
            when "01" & x"b75" => data <= x"0f";
            when "01" & x"b76" => data <= x"85";
            when "01" & x"b77" => data <= x"c8";
            when "01" & x"b78" => data <= x"b9";
            when "01" & x"b79" => data <= x"0e";
            when "01" & x"b7a" => data <= x"0f";
            when "01" & x"b7b" => data <= x"29";
            when "01" & x"b7c" => data <= x"03";
            when "01" & x"b7d" => data <= x"85";
            when "01" & x"b7e" => data <= x"c9";
            when "01" & x"b7f" => data <= x"c5";
            when "01" & x"b80" => data <= x"cb";
            when "01" & x"b81" => data <= x"d0";
            when "01" & x"b82" => data <= x"14";
            when "01" & x"b83" => data <= x"a5";
            when "01" & x"b84" => data <= x"c8";
            when "01" & x"b85" => data <= x"c5";
            when "01" & x"b86" => data <= x"ca";
            when "01" & x"b87" => data <= x"d0";
            when "01" & x"b88" => data <= x"0e";
            when "01" & x"b89" => data <= x"18";
            when "01" & x"b8a" => data <= x"65";
            when "01" & x"b8b" => data <= x"c6";
            when "01" & x"b8c" => data <= x"85";
            when "01" & x"b8d" => data <= x"ca";
            when "01" & x"b8e" => data <= x"a5";
            when "01" & x"b8f" => data <= x"cb";
            when "01" & x"b90" => data <= x"65";
            when "01" & x"b91" => data <= x"c7";
            when "01" & x"b92" => data <= x"85";
            when "01" & x"b93" => data <= x"cb";
            when "01" & x"b94" => data <= x"4c";
            when "01" & x"b95" => data <= x"b5";
            when "01" & x"b96" => data <= x"9b";
            when "01" & x"b97" => data <= x"a5";
            when "01" & x"b98" => data <= x"ca";
            when "01" & x"b99" => data <= x"99";
            when "01" & x"b9a" => data <= x"0f";
            when "01" & x"b9b" => data <= x"0f";
            when "01" & x"b9c" => data <= x"b9";
            when "01" & x"b9d" => data <= x"0e";
            when "01" & x"b9e" => data <= x"0f";
            when "01" & x"b9f" => data <= x"29";
            when "01" & x"ba0" => data <= x"fc";
            when "01" & x"ba1" => data <= x"05";
            when "01" & x"ba2" => data <= x"cb";
            when "01" & x"ba3" => data <= x"99";
            when "01" & x"ba4" => data <= x"0e";
            when "01" & x"ba5" => data <= x"0f";
            when "01" & x"ba6" => data <= x"a9";
            when "01" & x"ba7" => data <= x"00";
            when "01" & x"ba8" => data <= x"85";
            when "01" & x"ba9" => data <= x"a8";
            when "01" & x"baa" => data <= x"85";
            when "01" & x"bab" => data <= x"a9";
            when "01" & x"bac" => data <= x"20";
            when "01" & x"bad" => data <= x"b4";
            when "01" & x"bae" => data <= x"8a";
            when "01" & x"baf" => data <= x"20";
            when "01" & x"bb0" => data <= x"06";
            when "01" & x"bb1" => data <= x"9e";
            when "01" & x"bb2" => data <= x"20";
            when "01" & x"bb3" => data <= x"47";
            when "01" & x"bb4" => data <= x"83";
            when "01" & x"bb5" => data <= x"a4";
            when "01" & x"bb6" => data <= x"cc";
            when "01" & x"bb7" => data <= x"20";
            when "01" & x"bb8" => data <= x"01";
            when "01" & x"bb9" => data <= x"83";
            when "01" & x"bba" => data <= x"4c";
            when "01" & x"bbb" => data <= x"fb";
            when "01" & x"bbc" => data <= x"9a";
            when "01" & x"bbd" => data <= x"2c";
            when "01" & x"bbe" => data <= x"c8";
            when "01" & x"bbf" => data <= x"10";
            when "01" & x"bc0" => data <= x"10";
            when "01" & x"bc1" => data <= x"75";
            when "01" & x"bc2" => data <= x"20";
            when "01" & x"bc3" => data <= x"33";
            when "01" & x"bc4" => data <= x"80";
            when "01" & x"bc5" => data <= x"bd";
            when "01" & x"bc6" => data <= x"4e";
            when "01" & x"bc7" => data <= x"6f";
            when "01" & x"bc8" => data <= x"74";
            when "01" & x"bc9" => data <= x"20";
            when "01" & x"bca" => data <= x"65";
            when "01" & x"bcb" => data <= x"6e";
            when "01" & x"bcc" => data <= x"61";
            when "01" & x"bcd" => data <= x"62";
            when "01" & x"bce" => data <= x"6c";
            when "01" & x"bcf" => data <= x"65";
            when "01" & x"bd0" => data <= x"64";
            when "01" & x"bd1" => data <= x"00";
            when "01" & x"bd2" => data <= x"20";
            when "01" & x"bd3" => data <= x"bf";
            when "01" & x"bd4" => data <= x"86";
            when "01" & x"bd5" => data <= x"d0";
            when "01" & x"bd6" => data <= x"03";
            when "01" & x"bd7" => data <= x"4c";
            when "01" & x"bd8" => data <= x"06";
            when "01" & x"bd9" => data <= x"9a";
            when "01" & x"bda" => data <= x"20";
            when "01" & x"bdb" => data <= x"5d";
            when "01" & x"bdc" => data <= x"83";
            when "01" & x"bdd" => data <= x"8d";
            when "01" & x"bde" => data <= x"d2";
            when "01" & x"bdf" => data <= x"10";
            when "01" & x"be0" => data <= x"20";
            when "01" & x"be1" => data <= x"bf";
            when "01" & x"be2" => data <= x"86";
            when "01" & x"be3" => data <= x"f0";
            when "01" & x"be4" => data <= x"f2";
            when "01" & x"be5" => data <= x"20";
            when "01" & x"be6" => data <= x"5d";
            when "01" & x"be7" => data <= x"83";
            when "01" & x"be8" => data <= x"8d";
            when "01" & x"be9" => data <= x"d3";
            when "01" & x"bea" => data <= x"10";
            when "01" & x"beb" => data <= x"98";
            when "01" & x"bec" => data <= x"48";
            when "01" & x"bed" => data <= x"a9";
            when "01" & x"bee" => data <= x"00";
            when "01" & x"bef" => data <= x"85";
            when "01" & x"bf0" => data <= x"a9";
            when "01" & x"bf1" => data <= x"ad";
            when "01" & x"bf2" => data <= x"d3";
            when "01" & x"bf3" => data <= x"10";
            when "01" & x"bf4" => data <= x"cd";
            when "01" & x"bf5" => data <= x"d2";
            when "01" & x"bf6" => data <= x"10";
            when "01" & x"bf7" => data <= x"d0";
            when "01" & x"bf8" => data <= x"06";
            when "01" & x"bf9" => data <= x"a9";
            when "01" & x"bfa" => data <= x"ff";
            when "01" & x"bfb" => data <= x"85";
            when "01" & x"bfc" => data <= x"a9";
            when "01" & x"bfd" => data <= x"85";
            when "01" & x"bfe" => data <= x"aa";
            when "01" & x"bff" => data <= x"20";
            when "01" & x"c00" => data <= x"79";
            when "01" & x"c01" => data <= x"98";
            when "01" & x"c02" => data <= x"20";
            when "01" & x"c03" => data <= x"65";
            when "01" & x"c04" => data <= x"80";
            when "01" & x"c05" => data <= x"43";
            when "01" & x"c06" => data <= x"6f";
            when "01" & x"c07" => data <= x"70";
            when "01" & x"c08" => data <= x"79";
            when "01" & x"c09" => data <= x"69";
            when "01" & x"c0a" => data <= x"6e";
            when "01" & x"c0b" => data <= x"67";
            when "01" & x"c0c" => data <= x"20";
            when "01" & x"c0d" => data <= x"66";
            when "01" & x"c0e" => data <= x"72";
            when "01" & x"c0f" => data <= x"6f";
            when "01" & x"c10" => data <= x"6d";
            when "01" & x"c11" => data <= x"20";
            when "01" & x"c12" => data <= x"64";
            when "01" & x"c13" => data <= x"72";
            when "01" & x"c14" => data <= x"69";
            when "01" & x"c15" => data <= x"76";
            when "01" & x"c16" => data <= x"65";
            when "01" & x"c17" => data <= x"20";
            when "01" & x"c18" => data <= x"ad";
            when "01" & x"c19" => data <= x"d2";
            when "01" & x"c1a" => data <= x"10";
            when "01" & x"c1b" => data <= x"20";
            when "01" & x"c1c" => data <= x"ca";
            when "01" & x"c1d" => data <= x"80";
            when "01" & x"c1e" => data <= x"20";
            when "01" & x"c1f" => data <= x"65";
            when "01" & x"c20" => data <= x"80";
            when "01" & x"c21" => data <= x"20";
            when "01" & x"c22" => data <= x"74";
            when "01" & x"c23" => data <= x"6f";
            when "01" & x"c24" => data <= x"20";
            when "01" & x"c25" => data <= x"64";
            when "01" & x"c26" => data <= x"72";
            when "01" & x"c27" => data <= x"69";
            when "01" & x"c28" => data <= x"76";
            when "01" & x"c29" => data <= x"65";
            when "01" & x"c2a" => data <= x"20";
            when "01" & x"c2b" => data <= x"ad";
            when "01" & x"c2c" => data <= x"d3";
            when "01" & x"c2d" => data <= x"10";
            when "01" & x"c2e" => data <= x"20";
            when "01" & x"c2f" => data <= x"ca";
            when "01" & x"c30" => data <= x"80";
            when "01" & x"c31" => data <= x"20";
            when "01" & x"c32" => data <= x"9a";
            when "01" & x"c33" => data <= x"9f";
            when "01" & x"c34" => data <= x"68";
            when "01" & x"c35" => data <= x"a8";
            when "01" & x"c36" => data <= x"18";
            when "01" & x"c37" => data <= x"60";
            when "01" & x"c38" => data <= x"20";
            when "01" & x"c39" => data <= x"e1";
            when "01" & x"c3a" => data <= x"83";
            when "01" & x"c3b" => data <= x"24";
            when "01" & x"c3c" => data <= x"a9";
            when "01" & x"c3d" => data <= x"10";
            when "01" & x"c3e" => data <= x"0b";
            when "01" & x"c3f" => data <= x"a9";
            when "01" & x"c40" => data <= x"00";
            when "01" & x"c41" => data <= x"f0";
            when "01" & x"c42" => data <= x"0a";
            when "01" & x"c43" => data <= x"20";
            when "01" & x"c44" => data <= x"e1";
            when "01" & x"c45" => data <= x"83";
            when "01" & x"c46" => data <= x"24";
            when "01" & x"c47" => data <= x"a9";
            when "01" & x"c48" => data <= x"30";
            when "01" & x"c49" => data <= x"01";
            when "01" & x"c4a" => data <= x"60";
            when "01" & x"c4b" => data <= x"a9";
            when "01" & x"c4c" => data <= x"80";
            when "01" & x"c4d" => data <= x"c5";
            when "01" & x"c4e" => data <= x"aa";
            when "01" & x"c4f" => data <= x"f0";
            when "01" & x"c50" => data <= x"f9";
            when "01" & x"c51" => data <= x"85";
            when "01" & x"c52" => data <= x"aa";
            when "01" & x"c53" => data <= x"20";
            when "01" & x"c54" => data <= x"65";
            when "01" & x"c55" => data <= x"80";
            when "01" & x"c56" => data <= x"49";
            when "01" & x"c57" => data <= x"6e";
            when "01" & x"c58" => data <= x"73";
            when "01" & x"c59" => data <= x"65";
            when "01" & x"c5a" => data <= x"72";
            when "01" & x"c5b" => data <= x"74";
            when "01" & x"c5c" => data <= x"20";
            when "01" & x"c5d" => data <= x"ea";
            when "01" & x"c5e" => data <= x"24";
            when "01" & x"c5f" => data <= x"aa";
            when "01" & x"c60" => data <= x"30";
            when "01" & x"c61" => data <= x"0b";
            when "01" & x"c62" => data <= x"20";
            when "01" & x"c63" => data <= x"65";
            when "01" & x"c64" => data <= x"80";
            when "01" & x"c65" => data <= x"73";
            when "01" & x"c66" => data <= x"6f";
            when "01" & x"c67" => data <= x"75";
            when "01" & x"c68" => data <= x"72";
            when "01" & x"c69" => data <= x"63";
            when "01" & x"c6a" => data <= x"65";
            when "01" & x"c6b" => data <= x"90";
            when "01" & x"c6c" => data <= x"0f";
            when "01" & x"c6d" => data <= x"20";
            when "01" & x"c6e" => data <= x"65";
            when "01" & x"c6f" => data <= x"80";
            when "01" & x"c70" => data <= x"64";
            when "01" & x"c71" => data <= x"65";
            when "01" & x"c72" => data <= x"73";
            when "01" & x"c73" => data <= x"74";
            when "01" & x"c74" => data <= x"69";
            when "01" & x"c75" => data <= x"6e";
            when "01" & x"c76" => data <= x"61";
            when "01" & x"c77" => data <= x"74";
            when "01" & x"c78" => data <= x"69";
            when "01" & x"c79" => data <= x"6f";
            when "01" & x"c7a" => data <= x"6e";
            when "01" & x"c7b" => data <= x"ea";
            when "01" & x"c7c" => data <= x"20";
            when "01" & x"c7d" => data <= x"65";
            when "01" & x"c7e" => data <= x"80";
            when "01" & x"c7f" => data <= x"20";
            when "01" & x"c80" => data <= x"64";
            when "01" & x"c81" => data <= x"69";
            when "01" & x"c82" => data <= x"73";
            when "01" & x"c83" => data <= x"6b";
            when "01" & x"c84" => data <= x"20";
            when "01" & x"c85" => data <= x"61";
            when "01" & x"c86" => data <= x"6e";
            when "01" & x"c87" => data <= x"64";
            when "01" & x"c88" => data <= x"20";
            when "01" & x"c89" => data <= x"68";
            when "01" & x"c8a" => data <= x"69";
            when "01" & x"c8b" => data <= x"74";
            when "01" & x"c8c" => data <= x"20";
            when "01" & x"c8d" => data <= x"61";
            when "01" & x"c8e" => data <= x"20";
            when "01" & x"c8f" => data <= x"6b";
            when "01" & x"c90" => data <= x"65";
            when "01" & x"c91" => data <= x"79";
            when "01" & x"c92" => data <= x"ea";
            when "01" & x"c93" => data <= x"20";
            when "01" & x"c94" => data <= x"06";
            when "01" & x"c95" => data <= x"99";
            when "01" & x"c96" => data <= x"20";
            when "01" & x"c97" => data <= x"e0";
            when "01" & x"c98" => data <= x"ff";
            when "01" & x"c99" => data <= x"b0";
            when "01" & x"c9a" => data <= x"19";
            when "01" & x"c9b" => data <= x"4c";
            when "01" & x"c9c" => data <= x"9a";
            when "01" & x"c9d" => data <= x"9f";
            when "01" & x"c9e" => data <= x"20";
            when "01" & x"c9f" => data <= x"06";
            when "01" & x"ca0" => data <= x"99";
            when "01" & x"ca1" => data <= x"20";
            when "01" & x"ca2" => data <= x"e0";
            when "01" & x"ca3" => data <= x"ff";
            when "01" & x"ca4" => data <= x"b0";
            when "01" & x"ca5" => data <= x"0e";
            when "01" & x"ca6" => data <= x"29";
            when "01" & x"ca7" => data <= x"5f";
            when "01" & x"ca8" => data <= x"c9";
            when "01" & x"ca9" => data <= x"59";
            when "01" & x"caa" => data <= x"08";
            when "01" & x"cab" => data <= x"f0";
            when "01" & x"cac" => data <= x"02";
            when "01" & x"cad" => data <= x"a9";
            when "01" & x"cae" => data <= x"4e";
            when "01" & x"caf" => data <= x"20";
            when "01" & x"cb0" => data <= x"9c";
            when "01" & x"cb1" => data <= x"80";
            when "01" & x"cb2" => data <= x"28";
            when "01" & x"cb3" => data <= x"60";
            when "01" & x"cb4" => data <= x"a6";
            when "01" & x"cb5" => data <= x"b6";
            when "01" & x"cb6" => data <= x"9a";
            when "01" & x"cb7" => data <= x"60";
            when "01" & x"cb8" => data <= x"4c";
            when "01" & x"cb9" => data <= x"58";
            when "01" & x"cba" => data <= x"89";
            when "01" & x"cbb" => data <= x"20";
            when "01" & x"cbc" => data <= x"bd";
            when "01" & x"cbd" => data <= x"9b";
            when "01" & x"cbe" => data <= x"20";
            when "01" & x"cbf" => data <= x"d2";
            when "01" & x"cc0" => data <= x"9b";
            when "01" & x"cc1" => data <= x"a9";
            when "01" & x"cc2" => data <= x"00";
            when "01" & x"cc3" => data <= x"85";
            when "01" & x"cc4" => data <= x"c9";
            when "01" & x"cc5" => data <= x"85";
            when "01" & x"cc6" => data <= x"cb";
            when "01" & x"cc7" => data <= x"85";
            when "01" & x"cc8" => data <= x"ca";
            when "01" & x"cc9" => data <= x"85";
            when "01" & x"cca" => data <= x"c8";
            when "01" & x"ccb" => data <= x"85";
            when "01" & x"ccc" => data <= x"a8";
            when "01" & x"ccd" => data <= x"20";
            when "01" & x"cce" => data <= x"38";
            when "01" & x"ccf" => data <= x"9c";
            when "01" & x"cd0" => data <= x"ad";
            when "01" & x"cd1" => data <= x"d2";
            when "01" & x"cd2" => data <= x"10";
            when "01" & x"cd3" => data <= x"85";
            when "01" & x"cd4" => data <= x"cf";
            when "01" & x"cd5" => data <= x"20";
            when "01" & x"cd6" => data <= x"41";
            when "01" & x"cd7" => data <= x"af";
            when "01" & x"cd8" => data <= x"ad";
            when "01" & x"cd9" => data <= x"07";
            when "01" & x"cda" => data <= x"0f";
            when "01" & x"cdb" => data <= x"85";
            when "01" & x"cdc" => data <= x"c6";
            when "01" & x"cdd" => data <= x"ad";
            when "01" & x"cde" => data <= x"06";
            when "01" & x"cdf" => data <= x"0f";
            when "01" & x"ce0" => data <= x"29";
            when "01" & x"ce1" => data <= x"03";
            when "01" & x"ce2" => data <= x"85";
            when "01" & x"ce3" => data <= x"c7";
            when "01" & x"ce4" => data <= x"ad";
            when "01" & x"ce5" => data <= x"06";
            when "01" & x"ce6" => data <= x"0f";
            when "01" & x"ce7" => data <= x"29";
            when "01" & x"ce8" => data <= x"f0";
            when "01" & x"ce9" => data <= x"8d";
            when "01" & x"cea" => data <= x"d8";
            when "01" & x"ceb" => data <= x"10";
            when "01" & x"cec" => data <= x"20";
            when "01" & x"ced" => data <= x"43";
            when "01" & x"cee" => data <= x"9c";
            when "01" & x"cef" => data <= x"ad";
            when "01" & x"cf0" => data <= x"d3";
            when "01" & x"cf1" => data <= x"10";
            when "01" & x"cf2" => data <= x"85";
            when "01" & x"cf3" => data <= x"cf";
            when "01" & x"cf4" => data <= x"20";
            when "01" & x"cf5" => data <= x"41";
            when "01" & x"cf6" => data <= x"af";
            when "01" & x"cf7" => data <= x"ad";
            when "01" & x"cf8" => data <= x"06";
            when "01" & x"cf9" => data <= x"0f";
            when "01" & x"cfa" => data <= x"29";
            when "01" & x"cfb" => data <= x"03";
            when "01" & x"cfc" => data <= x"c5";
            when "01" & x"cfd" => data <= x"c7";
            when "01" & x"cfe" => data <= x"90";
            when "01" & x"cff" => data <= x"b8";
            when "01" & x"d00" => data <= x"d0";
            when "01" & x"d01" => data <= x"07";
            when "01" & x"d02" => data <= x"ad";
            when "01" & x"d03" => data <= x"07";
            when "01" & x"d04" => data <= x"0f";
            when "01" & x"d05" => data <= x"c5";
            when "01" & x"d06" => data <= x"c6";
            when "01" & x"d07" => data <= x"90";
            when "01" & x"d08" => data <= x"af";
            when "01" & x"d09" => data <= x"20";
            when "01" & x"d0a" => data <= x"06";
            when "01" & x"d0b" => data <= x"9e";
            when "01" & x"d0c" => data <= x"ad";
            when "01" & x"d0d" => data <= x"06";
            when "01" & x"d0e" => data <= x"0f";
            when "01" & x"d0f" => data <= x"48";
            when "01" & x"d10" => data <= x"ad";
            when "01" & x"d11" => data <= x"07";
            when "01" & x"d12" => data <= x"0f";
            when "01" & x"d13" => data <= x"48";
            when "01" & x"d14" => data <= x"20";
            when "01" & x"d15" => data <= x"41";
            when "01" & x"d16" => data <= x"af";
            when "01" & x"d17" => data <= x"68";
            when "01" & x"d18" => data <= x"8d";
            when "01" & x"d19" => data <= x"07";
            when "01" & x"d1a" => data <= x"0f";
            when "01" & x"d1b" => data <= x"68";
            when "01" & x"d1c" => data <= x"29";
            when "01" & x"d1d" => data <= x"0f";
            when "01" & x"d1e" => data <= x"0d";
            when "01" & x"d1f" => data <= x"d8";
            when "01" & x"d20" => data <= x"10";
            when "01" & x"d21" => data <= x"8d";
            when "01" & x"d22" => data <= x"06";
            when "01" & x"d23" => data <= x"0f";
            when "01" & x"d24" => data <= x"4c";
            when "01" & x"d25" => data <= x"b4";
            when "01" & x"d26" => data <= x"8a";
            when "01" & x"d27" => data <= x"20";
            when "01" & x"d28" => data <= x"5e";
            when "01" & x"d29" => data <= x"82";
            when "01" & x"d2a" => data <= x"20";
            when "01" & x"d2b" => data <= x"d2";
            when "01" & x"d2c" => data <= x"9b";
            when "01" & x"d2d" => data <= x"20";
            when "01" & x"d2e" => data <= x"bf";
            when "01" & x"d2f" => data <= x"86";
            when "01" & x"d30" => data <= x"d0";
            when "01" & x"d31" => data <= x"03";
            when "01" & x"d32" => data <= x"4c";
            when "01" & x"d33" => data <= x"06";
            when "01" & x"d34" => data <= x"9a";
            when "01" & x"d35" => data <= x"20";
            when "01" & x"d36" => data <= x"fe";
            when "01" & x"d37" => data <= x"80";
            when "01" & x"d38" => data <= x"20";
            when "01" & x"d39" => data <= x"38";
            when "01" & x"d3a" => data <= x"9c";
            when "01" & x"d3b" => data <= x"ad";
            when "01" & x"d3c" => data <= x"d2";
            when "01" & x"d3d" => data <= x"10";
            when "01" & x"d3e" => data <= x"20";
            when "01" & x"d3f" => data <= x"7e";
            when "01" & x"d40" => data <= x"87";
            when "01" & x"d41" => data <= x"20";
            when "01" & x"d42" => data <= x"96";
            when "01" & x"d43" => data <= x"82";
            when "01" & x"d44" => data <= x"b0";
            when "01" & x"d45" => data <= x"03";
            when "01" & x"d46" => data <= x"4c";
            when "01" & x"d47" => data <= x"76";
            when "01" & x"d48" => data <= x"82";
            when "01" & x"d49" => data <= x"84";
            when "01" & x"d4a" => data <= x"ab";
            when "01" & x"d4b" => data <= x"20";
            when "01" & x"d4c" => data <= x"01";
            when "01" & x"d4d" => data <= x"83";
            when "01" & x"d4e" => data <= x"a2";
            when "01" & x"d4f" => data <= x"00";
            when "01" & x"d50" => data <= x"b5";
            when "01" & x"d51" => data <= x"c7";
            when "01" & x"d52" => data <= x"9d";
            when "01" & x"d53" => data <= x"58";
            when "01" & x"d54" => data <= x"10";
            when "01" & x"d55" => data <= x"b9";
            when "01" & x"d56" => data <= x"08";
            when "01" & x"d57" => data <= x"0e";
            when "01" & x"d58" => data <= x"95";
            when "01" & x"d59" => data <= x"c7";
            when "01" & x"d5a" => data <= x"9d";
            when "01" & x"d5b" => data <= x"50";
            when "01" & x"d5c" => data <= x"10";
            when "01" & x"d5d" => data <= x"b9";
            when "01" & x"d5e" => data <= x"08";
            when "01" & x"d5f" => data <= x"0f";
            when "01" & x"d60" => data <= x"95";
            when "01" & x"d61" => data <= x"bd";
            when "01" & x"d62" => data <= x"9d";
            when "01" & x"d63" => data <= x"47";
            when "01" & x"d64" => data <= x"10";
            when "01" & x"d65" => data <= x"e8";
            when "01" & x"d66" => data <= x"c8";
            when "01" & x"d67" => data <= x"e0";
            when "01" & x"d68" => data <= x"08";
            when "01" & x"d69" => data <= x"d0";
            when "01" & x"d6a" => data <= x"e5";
            when "01" & x"d6b" => data <= x"a5";
            when "01" & x"d6c" => data <= x"c3";
            when "01" & x"d6d" => data <= x"20";
            when "01" & x"d6e" => data <= x"fd";
            when "01" & x"d6f" => data <= x"81";
            when "01" & x"d70" => data <= x"85";
            when "01" & x"d71" => data <= x"c5";
            when "01" & x"d72" => data <= x"a5";
            when "01" & x"d73" => data <= x"c1";
            when "01" & x"d74" => data <= x"18";
            when "01" & x"d75" => data <= x"69";
            when "01" & x"d76" => data <= x"ff";
            when "01" & x"d77" => data <= x"a5";
            when "01" & x"d78" => data <= x"c2";
            when "01" & x"d79" => data <= x"69";
            when "01" & x"d7a" => data <= x"00";
            when "01" & x"d7b" => data <= x"85";
            when "01" & x"d7c" => data <= x"c6";
            when "01" & x"d7d" => data <= x"a5";
            when "01" & x"d7e" => data <= x"c5";
            when "01" & x"d7f" => data <= x"69";
            when "01" & x"d80" => data <= x"00";
            when "01" & x"d81" => data <= x"85";
            when "01" & x"d82" => data <= x"c7";
            when "01" & x"d83" => data <= x"ad";
            when "01" & x"d84" => data <= x"4e";
            when "01" & x"d85" => data <= x"10";
            when "01" & x"d86" => data <= x"85";
            when "01" & x"d87" => data <= x"c8";
            when "01" & x"d88" => data <= x"ad";
            when "01" & x"d89" => data <= x"4d";
            when "01" & x"d8a" => data <= x"10";
            when "01" & x"d8b" => data <= x"29";
            when "01" & x"d8c" => data <= x"03";
            when "01" & x"d8d" => data <= x"85";
            when "01" & x"d8e" => data <= x"c9";
            when "01" & x"d8f" => data <= x"a9";
            when "01" & x"d90" => data <= x"ff";
            when "01" & x"d91" => data <= x"85";
            when "01" & x"d92" => data <= x"a8";
            when "01" & x"d93" => data <= x"20";
            when "01" & x"d94" => data <= x"06";
            when "01" & x"d95" => data <= x"9e";
            when "01" & x"d96" => data <= x"20";
            when "01" & x"d97" => data <= x"38";
            when "01" & x"d98" => data <= x"9c";
            when "01" & x"d99" => data <= x"ad";
            when "01" & x"d9a" => data <= x"d2";
            when "01" & x"d9b" => data <= x"10";
            when "01" & x"d9c" => data <= x"20";
            when "01" & x"d9d" => data <= x"7e";
            when "01" & x"d9e" => data <= x"87";
            when "01" & x"d9f" => data <= x"20";
            when "01" & x"da0" => data <= x"47";
            when "01" & x"da1" => data <= x"83";
            when "01" & x"da2" => data <= x"a2";
            when "01" & x"da3" => data <= x"07";
            when "01" & x"da4" => data <= x"bd";
            when "01" & x"da5" => data <= x"58";
            when "01" & x"da6" => data <= x"10";
            when "01" & x"da7" => data <= x"95";
            when "01" & x"da8" => data <= x"c7";
            when "01" & x"da9" => data <= x"ca";
            when "01" & x"daa" => data <= x"10";
            when "01" & x"dab" => data <= x"f8";
            when "01" & x"dac" => data <= x"a4";
            when "01" & x"dad" => data <= x"ab";
            when "01" & x"dae" => data <= x"8c";
            when "01" & x"daf" => data <= x"ce";
            when "01" & x"db0" => data <= x"10";
            when "01" & x"db1" => data <= x"20";
            when "01" & x"db2" => data <= x"9d";
            when "01" & x"db3" => data <= x"82";
            when "01" & x"db4" => data <= x"b0";
            when "01" & x"db5" => data <= x"93";
            when "01" & x"db6" => data <= x"60";
            when "01" & x"db7" => data <= x"20";
            when "01" & x"db8" => data <= x"f5";
            when "01" & x"db9" => data <= x"9d";
            when "01" & x"dba" => data <= x"20";
            when "01" & x"dbb" => data <= x"43";
            when "01" & x"dbc" => data <= x"9c";
            when "01" & x"dbd" => data <= x"ad";
            when "01" & x"dbe" => data <= x"d3";
            when "01" & x"dbf" => data <= x"10";
            when "01" & x"dc0" => data <= x"85";
            when "01" & x"dc1" => data <= x"cf";
            when "01" & x"dc2" => data <= x"a5";
            when "01" & x"dc3" => data <= x"ce";
            when "01" & x"dc4" => data <= x"48";
            when "01" & x"dc5" => data <= x"20";
            when "01" & x"dc6" => data <= x"47";
            when "01" & x"dc7" => data <= x"83";
            when "01" & x"dc8" => data <= x"20";
            when "01" & x"dc9" => data <= x"96";
            when "01" & x"dca" => data <= x"82";
            when "01" & x"dcb" => data <= x"90";
            when "01" & x"dcc" => data <= x"03";
            when "01" & x"dcd" => data <= x"20";
            when "01" & x"dce" => data <= x"d1";
            when "01" & x"dcf" => data <= x"82";
            when "01" & x"dd0" => data <= x"68";
            when "01" & x"dd1" => data <= x"85";
            when "01" & x"dd2" => data <= x"ce";
            when "01" & x"dd3" => data <= x"20";
            when "01" & x"dd4" => data <= x"3f";
            when "01" & x"dd5" => data <= x"8a";
            when "01" & x"dd6" => data <= x"20";
            when "01" & x"dd7" => data <= x"56";
            when "01" & x"dd8" => data <= x"8a";
            when "01" & x"dd9" => data <= x"a5";
            when "01" & x"dda" => data <= x"c4";
            when "01" & x"ddb" => data <= x"20";
            when "01" & x"ddc" => data <= x"fd";
            when "01" & x"ddd" => data <= x"81";
            when "01" & x"dde" => data <= x"85";
            when "01" & x"ddf" => data <= x"c6";
            when "01" & x"de0" => data <= x"20";
            when "01" & x"de1" => data <= x"9d";
            when "01" & x"de2" => data <= x"89";
            when "01" & x"de3" => data <= x"a5";
            when "01" & x"de4" => data <= x"c4";
            when "01" & x"de5" => data <= x"29";
            when "01" & x"de6" => data <= x"03";
            when "01" & x"de7" => data <= x"48";
            when "01" & x"de8" => data <= x"a5";
            when "01" & x"de9" => data <= x"c5";
            when "01" & x"dea" => data <= x"48";
            when "01" & x"deb" => data <= x"20";
            when "01" & x"dec" => data <= x"f5";
            when "01" & x"ded" => data <= x"9d";
            when "01" & x"dee" => data <= x"68";
            when "01" & x"def" => data <= x"85";
            when "01" & x"df0" => data <= x"ca";
            when "01" & x"df1" => data <= x"68";
            when "01" & x"df2" => data <= x"85";
            when "01" & x"df3" => data <= x"cb";
            when "01" & x"df4" => data <= x"60";
            when "01" & x"df5" => data <= x"a2";
            when "01" & x"df6" => data <= x"11";
            when "01" & x"df7" => data <= x"bd";
            when "01" & x"df8" => data <= x"45";
            when "01" & x"df9" => data <= x"10";
            when "01" & x"dfa" => data <= x"b4";
            when "01" & x"dfb" => data <= x"bc";
            when "01" & x"dfc" => data <= x"95";
            when "01" & x"dfd" => data <= x"bc";
            when "01" & x"dfe" => data <= x"98";
            when "01" & x"dff" => data <= x"9d";
            when "01" & x"e00" => data <= x"45";
            when "01" & x"e01" => data <= x"10";
            when "01" & x"e02" => data <= x"ca";
            when "01" & x"e03" => data <= x"10";
            when "01" & x"e04" => data <= x"f2";
            when "01" & x"e05" => data <= x"60";
            when "01" & x"e06" => data <= x"20";
            when "01" & x"e07" => data <= x"8d";
            when "01" & x"e08" => data <= x"a0";
            when "01" & x"e09" => data <= x"a9";
            when "01" & x"e0a" => data <= x"00";
            when "01" & x"e0b" => data <= x"85";
            when "01" & x"e0c" => data <= x"be";
            when "01" & x"e0d" => data <= x"85";
            when "01" & x"e0e" => data <= x"c2";
            when "01" & x"e0f" => data <= x"a5";
            when "01" & x"e10" => data <= x"c6";
            when "01" & x"e11" => data <= x"a8";
            when "01" & x"e12" => data <= x"cd";
            when "01" & x"e13" => data <= x"d1";
            when "01" & x"e14" => data <= x"10";
            when "01" & x"e15" => data <= x"a5";
            when "01" & x"e16" => data <= x"c7";
            when "01" & x"e17" => data <= x"e9";
            when "01" & x"e18" => data <= x"00";
            when "01" & x"e19" => data <= x"90";
            when "01" & x"e1a" => data <= x"03";
            when "01" & x"e1b" => data <= x"ac";
            when "01" & x"e1c" => data <= x"d1";
            when "01" & x"e1d" => data <= x"10";
            when "01" & x"e1e" => data <= x"84";
            when "01" & x"e1f" => data <= x"c3";
            when "01" & x"e20" => data <= x"a5";
            when "01" & x"e21" => data <= x"c8";
            when "01" & x"e22" => data <= x"85";
            when "01" & x"e23" => data <= x"c5";
            when "01" & x"e24" => data <= x"a5";
            when "01" & x"e25" => data <= x"c9";
            when "01" & x"e26" => data <= x"85";
            when "01" & x"e27" => data <= x"c4";
            when "01" & x"e28" => data <= x"ad";
            when "01" & x"e29" => data <= x"d0";
            when "01" & x"e2a" => data <= x"10";
            when "01" & x"e2b" => data <= x"85";
            when "01" & x"e2c" => data <= x"bf";
            when "01" & x"e2d" => data <= x"ad";
            when "01" & x"e2e" => data <= x"d2";
            when "01" & x"e2f" => data <= x"10";
            when "01" & x"e30" => data <= x"85";
            when "01" & x"e31" => data <= x"cf";
            when "01" & x"e32" => data <= x"20";
            when "01" & x"e33" => data <= x"38";
            when "01" & x"e34" => data <= x"9c";
            when "01" & x"e35" => data <= x"20";
            when "01" & x"e36" => data <= x"3e";
            when "01" & x"e37" => data <= x"be";
            when "01" & x"e38" => data <= x"20";
            when "01" & x"e39" => data <= x"c6";
            when "01" & x"e3a" => data <= x"87";
            when "01" & x"e3b" => data <= x"ad";
            when "01" & x"e3c" => data <= x"d3";
            when "01" & x"e3d" => data <= x"10";
            when "01" & x"e3e" => data <= x"85";
            when "01" & x"e3f" => data <= x"cf";
            when "01" & x"e40" => data <= x"24";
            when "01" & x"e41" => data <= x"a8";
            when "01" & x"e42" => data <= x"10";
            when "01" & x"e43" => data <= x"07";
            when "01" & x"e44" => data <= x"20";
            when "01" & x"e45" => data <= x"b7";
            when "01" & x"e46" => data <= x"9d";
            when "01" & x"e47" => data <= x"a9";
            when "01" & x"e48" => data <= x"00";
            when "01" & x"e49" => data <= x"85";
            when "01" & x"e4a" => data <= x"a8";
            when "01" & x"e4b" => data <= x"a5";
            when "01" & x"e4c" => data <= x"ca";
            when "01" & x"e4d" => data <= x"85";
            when "01" & x"e4e" => data <= x"c5";
            when "01" & x"e4f" => data <= x"a5";
            when "01" & x"e50" => data <= x"cb";
            when "01" & x"e51" => data <= x"85";
            when "01" & x"e52" => data <= x"c4";
            when "01" & x"e53" => data <= x"ad";
            when "01" & x"e54" => data <= x"d0";
            when "01" & x"e55" => data <= x"10";
            when "01" & x"e56" => data <= x"85";
            when "01" & x"e57" => data <= x"bf";
            when "01" & x"e58" => data <= x"20";
            when "01" & x"e59" => data <= x"43";
            when "01" & x"e5a" => data <= x"9c";
            when "01" & x"e5b" => data <= x"20";
            when "01" & x"e5c" => data <= x"3e";
            when "01" & x"e5d" => data <= x"be";
            when "01" & x"e5e" => data <= x"20";
            when "01" & x"e5f" => data <= x"8f";
            when "01" & x"e60" => data <= x"87";
            when "01" & x"e61" => data <= x"a5";
            when "01" & x"e62" => data <= x"c3";
            when "01" & x"e63" => data <= x"18";
            when "01" & x"e64" => data <= x"65";
            when "01" & x"e65" => data <= x"ca";
            when "01" & x"e66" => data <= x"85";
            when "01" & x"e67" => data <= x"ca";
            when "01" & x"e68" => data <= x"90";
            when "01" & x"e69" => data <= x"02";
            when "01" & x"e6a" => data <= x"e6";
            when "01" & x"e6b" => data <= x"cb";
            when "01" & x"e6c" => data <= x"a5";
            when "01" & x"e6d" => data <= x"c3";
            when "01" & x"e6e" => data <= x"18";
            when "01" & x"e6f" => data <= x"65";
            when "01" & x"e70" => data <= x"c8";
            when "01" & x"e71" => data <= x"85";
            when "01" & x"e72" => data <= x"c8";
            when "01" & x"e73" => data <= x"90";
            when "01" & x"e74" => data <= x"02";
            when "01" & x"e75" => data <= x"e6";
            when "01" & x"e76" => data <= x"c9";
            when "01" & x"e77" => data <= x"38";
            when "01" & x"e78" => data <= x"a5";
            when "01" & x"e79" => data <= x"c6";
            when "01" & x"e7a" => data <= x"e5";
            when "01" & x"e7b" => data <= x"c3";
            when "01" & x"e7c" => data <= x"85";
            when "01" & x"e7d" => data <= x"c6";
            when "01" & x"e7e" => data <= x"b0";
            when "01" & x"e7f" => data <= x"02";
            when "01" & x"e80" => data <= x"c6";
            when "01" & x"e81" => data <= x"c7";
            when "01" & x"e82" => data <= x"05";
            when "01" & x"e83" => data <= x"c7";
            when "01" & x"e84" => data <= x"d0";
            when "01" & x"e85" => data <= x"89";
            when "01" & x"e86" => data <= x"60";
            when "01" & x"e87" => data <= x"20";
            when "01" & x"e88" => data <= x"d7";
            when "01" & x"e89" => data <= x"9f";
            when "01" & x"e8a" => data <= x"a9";
            when "01" & x"e8b" => data <= x"00";
            when "01" & x"e8c" => data <= x"f0";
            when "01" & x"e8d" => data <= x"05";
            when "01" & x"e8e" => data <= x"20";
            when "01" & x"e8f" => data <= x"d7";
            when "01" & x"e90" => data <= x"9f";
            when "01" & x"e91" => data <= x"a9";
            when "01" & x"e92" => data <= x"ff";
            when "01" & x"e93" => data <= x"85";
            when "01" & x"e94" => data <= x"ab";
            when "01" & x"e95" => data <= x"a9";
            when "01" & x"e96" => data <= x"c0";
            when "01" & x"e97" => data <= x"20";
            when "01" & x"e98" => data <= x"ce";
            when "01" & x"e99" => data <= x"ff";
            when "01" & x"e9a" => data <= x"a8";
            when "01" & x"e9b" => data <= x"a9";
            when "01" & x"e9c" => data <= x"0d";
            when "01" & x"e9d" => data <= x"c0";
            when "01" & x"e9e" => data <= x"00";
            when "01" & x"e9f" => data <= x"d0";
            when "01" & x"ea0" => data <= x"1e";
            when "01" & x"ea1" => data <= x"4c";
            when "01" & x"ea2" => data <= x"76";
            when "01" & x"ea3" => data <= x"82";
            when "01" & x"ea4" => data <= x"20";
            when "01" & x"ea5" => data <= x"d7";
            when "01" & x"ea6" => data <= x"ff";
            when "01" & x"ea7" => data <= x"b0";
            when "01" & x"ea8" => data <= x"1e";
            when "01" & x"ea9" => data <= x"c9";
            when "01" & x"eaa" => data <= x"0a";
            when "01" & x"eab" => data <= x"f0";
            when "01" & x"eac" => data <= x"f7";
            when "01" & x"ead" => data <= x"28";
            when "01" & x"eae" => data <= x"d0";
            when "01" & x"eaf" => data <= x"08";
            when "01" & x"eb0" => data <= x"48";
            when "01" & x"eb1" => data <= x"20";
            when "01" & x"eb2" => data <= x"a2";
            when "01" & x"eb3" => data <= x"9f";
            when "01" & x"eb4" => data <= x"20";
            when "01" & x"eb5" => data <= x"ce";
            when "01" & x"eb6" => data <= x"9f";
            when "01" & x"eb7" => data <= x"68";
            when "01" & x"eb8" => data <= x"20";
            when "01" & x"eb9" => data <= x"e3";
            when "01" & x"eba" => data <= x"ff";
            when "01" & x"ebb" => data <= x"24";
            when "01" & x"ebc" => data <= x"ff";
            when "01" & x"ebd" => data <= x"30";
            when "01" & x"ebe" => data <= x"09";
            when "01" & x"ebf" => data <= x"25";
            when "01" & x"ec0" => data <= x"ab";
            when "01" & x"ec1" => data <= x"c9";
            when "01" & x"ec2" => data <= x"0d";
            when "01" & x"ec3" => data <= x"08";
            when "01" & x"ec4" => data <= x"4c";
            when "01" & x"ec5" => data <= x"a4";
            when "01" & x"ec6" => data <= x"9e";
            when "01" & x"ec7" => data <= x"28";
            when "01" & x"ec8" => data <= x"20";
            when "01" & x"ec9" => data <= x"9a";
            when "01" & x"eca" => data <= x"9f";
            when "01" & x"ecb" => data <= x"a9";
            when "01" & x"ecc" => data <= x"00";
            when "01" & x"ecd" => data <= x"4c";
            when "01" & x"ece" => data <= x"ce";
            when "01" & x"ecf" => data <= x"ff";
            when "01" & x"ed0" => data <= x"20";
            when "01" & x"ed1" => data <= x"d7";
            when "01" & x"ed2" => data <= x"9f";
            when "01" & x"ed3" => data <= x"a9";
            when "01" & x"ed4" => data <= x"c0";
            when "01" & x"ed5" => data <= x"20";
            when "01" & x"ed6" => data <= x"ce";
            when "01" & x"ed7" => data <= x"ff";
            when "01" & x"ed8" => data <= x"a8";
            when "01" & x"ed9" => data <= x"f0";
            when "01" & x"eda" => data <= x"c6";
            when "01" & x"edb" => data <= x"a6";
            when "01" & x"edc" => data <= x"f4";
            when "01" & x"edd" => data <= x"bd";
            when "01" & x"ede" => data <= x"f0";
            when "01" & x"edf" => data <= x"0d";
            when "01" & x"ee0" => data <= x"85";
            when "01" & x"ee1" => data <= x"ad";
            when "01" & x"ee2" => data <= x"e6";
            when "01" & x"ee3" => data <= x"ad";
            when "01" & x"ee4" => data <= x"24";
            when "01" & x"ee5" => data <= x"ff";
            when "01" & x"ee6" => data <= x"30";
            when "01" & x"ee7" => data <= x"e3";
            when "01" & x"ee8" => data <= x"a5";
            when "01" & x"ee9" => data <= x"a9";
            when "01" & x"eea" => data <= x"20";
            when "01" & x"eeb" => data <= x"c2";
            when "01" & x"eec" => data <= x"80";
            when "01" & x"eed" => data <= x"a5";
            when "01" & x"eee" => data <= x"a8";
            when "01" & x"eef" => data <= x"20";
            when "01" & x"ef0" => data <= x"c2";
            when "01" & x"ef1" => data <= x"80";
            when "01" & x"ef2" => data <= x"20";
            when "01" & x"ef3" => data <= x"ce";
            when "01" & x"ef4" => data <= x"9f";
            when "01" & x"ef5" => data <= x"a9";
            when "01" & x"ef6" => data <= x"07";
            when "01" & x"ef7" => data <= x"85";
            when "01" & x"ef8" => data <= x"ac";
            when "01" & x"ef9" => data <= x"a2";
            when "01" & x"efa" => data <= x"00";
            when "01" & x"efb" => data <= x"20";
            when "01" & x"efc" => data <= x"d7";
            when "01" & x"efd" => data <= x"ff";
            when "01" & x"efe" => data <= x"b0";
            when "01" & x"eff" => data <= x"0d";
            when "01" & x"f00" => data <= x"81";
            when "01" & x"f01" => data <= x"ac";
            when "01" & x"f02" => data <= x"20";
            when "01" & x"f03" => data <= x"c2";
            when "01" & x"f04" => data <= x"80";
            when "01" & x"f05" => data <= x"20";
            when "01" & x"f06" => data <= x"ce";
            when "01" & x"f07" => data <= x"9f";
            when "01" & x"f08" => data <= x"c6";
            when "01" & x"f09" => data <= x"ac";
            when "01" & x"f0a" => data <= x"10";
            when "01" & x"f0b" => data <= x"ef";
            when "01" & x"f0c" => data <= x"18";
            when "01" & x"f0d" => data <= x"08";
            when "01" & x"f0e" => data <= x"90";
            when "01" & x"f0f" => data <= x"0e";
            when "01" & x"f10" => data <= x"20";
            when "01" & x"f11" => data <= x"65";
            when "01" & x"f12" => data <= x"80";
            when "01" & x"f13" => data <= x"2a";
            when "01" & x"f14" => data <= x"2a";
            when "01" & x"f15" => data <= x"20";
            when "01" & x"f16" => data <= x"a9";
            when "01" & x"f17" => data <= x"00";
            when "01" & x"f18" => data <= x"81";
            when "01" & x"f19" => data <= x"ac";
            when "01" & x"f1a" => data <= x"c6";
            when "01" & x"f1b" => data <= x"ac";
            when "01" & x"f1c" => data <= x"10";
            when "01" & x"f1d" => data <= x"f2";
            when "01" & x"f1e" => data <= x"a9";
            when "01" & x"f1f" => data <= x"07";
            when "01" & x"f20" => data <= x"85";
            when "01" & x"f21" => data <= x"ac";
            when "01" & x"f22" => data <= x"a1";
            when "01" & x"f23" => data <= x"ac";
            when "01" & x"f24" => data <= x"c9";
            when "01" & x"f25" => data <= x"7f";
            when "01" & x"f26" => data <= x"b0";
            when "01" & x"f27" => data <= x"04";
            when "01" & x"f28" => data <= x"c9";
            when "01" & x"f29" => data <= x"20";
            when "01" & x"f2a" => data <= x"b0";
            when "01" & x"f2b" => data <= x"02";
            when "01" & x"f2c" => data <= x"a9";
            when "01" & x"f2d" => data <= x"2e";
            when "01" & x"f2e" => data <= x"20";
            when "01" & x"f2f" => data <= x"e3";
            when "01" & x"f30" => data <= x"ff";
            when "01" & x"f31" => data <= x"c6";
            when "01" & x"f32" => data <= x"ac";
            when "01" & x"f33" => data <= x"10";
            when "01" & x"f34" => data <= x"ed";
            when "01" & x"f35" => data <= x"20";
            when "01" & x"f36" => data <= x"9a";
            when "01" & x"f37" => data <= x"9f";
            when "01" & x"f38" => data <= x"a9";
            when "01" & x"f39" => data <= x"08";
            when "01" & x"f3a" => data <= x"18";
            when "01" & x"f3b" => data <= x"65";
            when "01" & x"f3c" => data <= x"a8";
            when "01" & x"f3d" => data <= x"85";
            when "01" & x"f3e" => data <= x"a8";
            when "01" & x"f3f" => data <= x"90";
            when "01" & x"f40" => data <= x"02";
            when "01" & x"f41" => data <= x"e6";
            when "01" & x"f42" => data <= x"a9";
            when "01" & x"f43" => data <= x"28";
            when "01" & x"f44" => data <= x"90";
            when "01" & x"f45" => data <= x"9e";
            when "01" & x"f46" => data <= x"b0";
            when "01" & x"f47" => data <= x"83";
            when "01" & x"f48" => data <= x"20";
            when "01" & x"f49" => data <= x"d7";
            when "01" & x"f4a" => data <= x"9f";
            when "01" & x"f4b" => data <= x"a9";
            when "01" & x"f4c" => data <= x"80";
            when "01" & x"f4d" => data <= x"20";
            when "01" & x"f4e" => data <= x"ce";
            when "01" & x"f4f" => data <= x"ff";
            when "01" & x"f50" => data <= x"85";
            when "01" & x"f51" => data <= x"ab";
            when "01" & x"f52" => data <= x"20";
            when "01" & x"f53" => data <= x"a2";
            when "01" & x"f54" => data <= x"9f";
            when "01" & x"f55" => data <= x"20";
            when "01" & x"f56" => data <= x"ce";
            when "01" & x"f57" => data <= x"9f";
            when "01" & x"f58" => data <= x"a6";
            when "01" & x"f59" => data <= x"f4";
            when "01" & x"f5a" => data <= x"bc";
            when "01" & x"f5b" => data <= x"f0";
            when "01" & x"f5c" => data <= x"0d";
            when "01" & x"f5d" => data <= x"c8";
            when "01" & x"f5e" => data <= x"84";
            when "01" & x"f5f" => data <= x"ad";
            when "01" & x"f60" => data <= x"a2";
            when "01" & x"f61" => data <= x"ac";
            when "01" & x"f62" => data <= x"a0";
            when "01" & x"f63" => data <= x"ff";
            when "01" & x"f64" => data <= x"84";
            when "01" & x"f65" => data <= x"ae";
            when "01" & x"f66" => data <= x"84";
            when "01" & x"f67" => data <= x"b0";
            when "01" & x"f68" => data <= x"c8";
            when "01" & x"f69" => data <= x"84";
            when "01" & x"f6a" => data <= x"ac";
            when "01" & x"f6b" => data <= x"84";
            when "01" & x"f6c" => data <= x"af";
            when "01" & x"f6d" => data <= x"98";
            when "01" & x"f6e" => data <= x"20";
            when "01" & x"f6f" => data <= x"f1";
            when "01" & x"f70" => data <= x"ff";
            when "01" & x"f71" => data <= x"08";
            when "01" & x"f72" => data <= x"84";
            when "01" & x"f73" => data <= x"aa";
            when "01" & x"f74" => data <= x"a4";
            when "01" & x"f75" => data <= x"ab";
            when "01" & x"f76" => data <= x"a2";
            when "01" & x"f77" => data <= x"00";
            when "01" & x"f78" => data <= x"f0";
            when "01" & x"f79" => data <= x"07";
            when "01" & x"f7a" => data <= x"a1";
            when "01" & x"f7b" => data <= x"ac";
            when "01" & x"f7c" => data <= x"20";
            when "01" & x"f7d" => data <= x"d4";
            when "01" & x"f7e" => data <= x"ff";
            when "01" & x"f7f" => data <= x"e6";
            when "01" & x"f80" => data <= x"ac";
            when "01" & x"f81" => data <= x"a5";
            when "01" & x"f82" => data <= x"ac";
            when "01" & x"f83" => data <= x"c5";
            when "01" & x"f84" => data <= x"aa";
            when "01" & x"f85" => data <= x"d0";
            when "01" & x"f86" => data <= x"f3";
            when "01" & x"f87" => data <= x"28";
            when "01" & x"f88" => data <= x"b0";
            when "01" & x"f89" => data <= x"08";
            when "01" & x"f8a" => data <= x"a9";
            when "01" & x"f8b" => data <= x"0d";
            when "01" & x"f8c" => data <= x"20";
            when "01" & x"f8d" => data <= x"d4";
            when "01" & x"f8e" => data <= x"ff";
            when "01" & x"f8f" => data <= x"4c";
            when "01" & x"f90" => data <= x"52";
            when "01" & x"f91" => data <= x"9f";
            when "01" & x"f92" => data <= x"a9";
            when "01" & x"f93" => data <= x"7e";
            when "01" & x"f94" => data <= x"20";
            when "01" & x"f95" => data <= x"f4";
            when "01" & x"f96" => data <= x"ff";
            when "01" & x"f97" => data <= x"20";
            when "01" & x"f98" => data <= x"cb";
            when "01" & x"f99" => data <= x"9e";
            when "01" & x"f9a" => data <= x"48";
            when "01" & x"f9b" => data <= x"a9";
            when "01" & x"f9c" => data <= x"0d";
            when "01" & x"f9d" => data <= x"20";
            when "01" & x"f9e" => data <= x"9c";
            when "01" & x"f9f" => data <= x"80";
            when "01" & x"fa0" => data <= x"68";
            when "01" & x"fa1" => data <= x"60";
            when "01" & x"fa2" => data <= x"f8";
            when "01" & x"fa3" => data <= x"18";
            when "01" & x"fa4" => data <= x"a5";
            when "01" & x"fa5" => data <= x"a8";
            when "01" & x"fa6" => data <= x"69";
            when "01" & x"fa7" => data <= x"01";
            when "01" & x"fa8" => data <= x"85";
            when "01" & x"fa9" => data <= x"a8";
            when "01" & x"faa" => data <= x"a5";
            when "01" & x"fab" => data <= x"a9";
            when "01" & x"fac" => data <= x"69";
            when "01" & x"fad" => data <= x"00";
            when "01" & x"fae" => data <= x"85";
            when "01" & x"faf" => data <= x"a9";
            when "01" & x"fb0" => data <= x"d8";
            when "01" & x"fb1" => data <= x"18";
            when "01" & x"fb2" => data <= x"20";
            when "01" & x"fb3" => data <= x"b7";
            when "01" & x"fb4" => data <= x"9f";
            when "01" & x"fb5" => data <= x"a5";
            when "01" & x"fb6" => data <= x"a8";
            when "01" & x"fb7" => data <= x"48";
            when "01" & x"fb8" => data <= x"08";
            when "01" & x"fb9" => data <= x"20";
            when "01" & x"fba" => data <= x"05";
            when "01" & x"fbb" => data <= x"82";
            when "01" & x"fbc" => data <= x"28";
            when "01" & x"fbd" => data <= x"20";
            when "01" & x"fbe" => data <= x"c1";
            when "01" & x"fbf" => data <= x"9f";
            when "01" & x"fc0" => data <= x"68";
            when "01" & x"fc1" => data <= x"aa";
            when "01" & x"fc2" => data <= x"b0";
            when "01" & x"fc3" => data <= x"02";
            when "01" & x"fc4" => data <= x"f0";
            when "01" & x"fc5" => data <= x"08";
            when "01" & x"fc6" => data <= x"20";
            when "01" & x"fc7" => data <= x"ca";
            when "01" & x"fc8" => data <= x"80";
            when "01" & x"fc9" => data <= x"38";
            when "01" & x"fca" => data <= x"60";
            when "01" & x"fcb" => data <= x"20";
            when "01" & x"fcc" => data <= x"ce";
            when "01" & x"fcd" => data <= x"9f";
            when "01" & x"fce" => data <= x"48";
            when "01" & x"fcf" => data <= x"a9";
            when "01" & x"fd0" => data <= x"20";
            when "01" & x"fd1" => data <= x"20";
            when "01" & x"fd2" => data <= x"9c";
            when "01" & x"fd3" => data <= x"80";
            when "01" & x"fd4" => data <= x"68";
            when "01" & x"fd5" => data <= x"18";
            when "01" & x"fd6" => data <= x"60";
            when "01" & x"fd7" => data <= x"ba";
            when "01" & x"fd8" => data <= x"a9";
            when "01" & x"fd9" => data <= x"00";
            when "01" & x"fda" => data <= x"9d";
            when "01" & x"fdb" => data <= x"07";
            when "01" & x"fdc" => data <= x"01";
            when "01" & x"fdd" => data <= x"88";
            when "01" & x"fde" => data <= x"c8";
            when "01" & x"fdf" => data <= x"b1";
            when "01" & x"fe0" => data <= x"f2";
            when "01" & x"fe1" => data <= x"c9";
            when "01" & x"fe2" => data <= x"20";
            when "01" & x"fe3" => data <= x"f0";
            when "01" & x"fe4" => data <= x"f9";
            when "01" & x"fe5" => data <= x"c9";
            when "01" & x"fe6" => data <= x"0d";
            when "01" & x"fe7" => data <= x"d0";
            when "01" & x"fe8" => data <= x"03";
            when "01" & x"fe9" => data <= x"4c";
            when "01" & x"fea" => data <= x"06";
            when "01" & x"feb" => data <= x"9a";
            when "01" & x"fec" => data <= x"a9";
            when "01" & x"fed" => data <= x"00";
            when "01" & x"fee" => data <= x"85";
            when "01" & x"fef" => data <= x"a8";
            when "01" & x"ff0" => data <= x"85";
            when "01" & x"ff1" => data <= x"a9";
            when "01" & x"ff2" => data <= x"48";
            when "01" & x"ff3" => data <= x"98";
            when "01" & x"ff4" => data <= x"18";
            when "01" & x"ff5" => data <= x"65";
            when "01" & x"ff6" => data <= x"f2";
            when "01" & x"ff7" => data <= x"aa";
            when "01" & x"ff8" => data <= x"a5";
            when "01" & x"ff9" => data <= x"f3";
            when "01" & x"ffa" => data <= x"69";
            when "01" & x"ffb" => data <= x"00";
            when "01" & x"ffc" => data <= x"a8";
            when "01" & x"ffd" => data <= x"68";
            when "01" & x"ffe" => data <= x"60";
            when "01" & x"fff" => data <= x"6d";
            when "10" & x"000" => data <= x"20";
            when "10" & x"001" => data <= x"80";
            when "10" & x"002" => data <= x"a1";
            when "10" & x"003" => data <= x"68";
            when "10" & x"004" => data <= x"85";
            when "10" & x"005" => data <= x"b8";
            when "10" & x"006" => data <= x"68";
            when "10" & x"007" => data <= x"85";
            when "10" & x"008" => data <= x"b9";
            when "10" & x"009" => data <= x"20";
            when "10" & x"00a" => data <= x"0f";
            when "10" & x"00b" => data <= x"a0";
            when "10" & x"00c" => data <= x"4c";
            when "10" & x"00d" => data <= x"00";
            when "10" & x"00e" => data <= x"01";
            when "10" & x"00f" => data <= x"a0";
            when "10" & x"010" => data <= x"00";
            when "10" & x"011" => data <= x"8c";
            when "10" & x"012" => data <= x"00";
            when "10" & x"013" => data <= x"01";
            when "10" & x"014" => data <= x"c8";
            when "10" & x"015" => data <= x"f0";
            when "10" & x"016" => data <= x"07";
            when "10" & x"017" => data <= x"b1";
            when "10" & x"018" => data <= x"b8";
            when "10" & x"019" => data <= x"99";
            when "10" & x"01a" => data <= x"00";
            when "10" & x"01b" => data <= x"01";
            when "10" & x"01c" => data <= x"d0";
            when "10" & x"01d" => data <= x"f6";
            when "10" & x"01e" => data <= x"60";
            when "10" & x"01f" => data <= x"a2";
            when "10" & x"020" => data <= x"ff";
            when "10" & x"021" => data <= x"d0";
            when "10" & x"022" => data <= x"02";
            when "10" & x"023" => data <= x"a2";
            when "10" & x"024" => data <= x"00";
            when "10" & x"025" => data <= x"a0";
            when "10" & x"026" => data <= x"ff";
            when "10" & x"027" => data <= x"8c";
            when "10" & x"028" => data <= x"82";
            when "10" & x"029" => data <= x"10";
            when "10" & x"02a" => data <= x"85";
            when "10" & x"02b" => data <= x"b0";
            when "10" & x"02c" => data <= x"86";
            when "10" & x"02d" => data <= x"b1";
            when "10" & x"02e" => data <= x"8d";
            when "10" & x"02f" => data <= x"02";
            when "10" & x"030" => data <= x"0d";
            when "10" & x"031" => data <= x"20";
            when "10" & x"032" => data <= x"80";
            when "10" & x"033" => data <= x"a1";
            when "10" & x"034" => data <= x"68";
            when "10" & x"035" => data <= x"85";
            when "10" & x"036" => data <= x"b8";
            when "10" & x"037" => data <= x"68";
            when "10" & x"038" => data <= x"85";
            when "10" & x"039" => data <= x"b9";
            when "10" & x"03a" => data <= x"20";
            when "10" & x"03b" => data <= x"0f";
            when "10" & x"03c" => data <= x"a0";
            when "10" & x"03d" => data <= x"a5";
            when "10" & x"03e" => data <= x"b0";
            when "10" & x"03f" => data <= x"20";
            when "10" & x"040" => data <= x"69";
            when "10" & x"041" => data <= x"a0";
            when "10" & x"042" => data <= x"a5";
            when "10" & x"043" => data <= x"b1";
            when "10" & x"044" => data <= x"f0";
            when "10" & x"045" => data <= x"1b";
            when "10" & x"046" => data <= x"a9";
            when "10" & x"047" => data <= x"2f";
            when "10" & x"048" => data <= x"99";
            when "10" & x"049" => data <= x"00";
            when "10" & x"04a" => data <= x"01";
            when "10" & x"04b" => data <= x"c8";
            when "10" & x"04c" => data <= x"ae";
            when "10" & x"04d" => data <= x"41";
            when "10" & x"04e" => data <= x"0d";
            when "10" & x"04f" => data <= x"bd";
            when "10" & x"050" => data <= x"44";
            when "10" & x"051" => data <= x"0d";
            when "10" & x"052" => data <= x"20";
            when "10" & x"053" => data <= x"69";
            when "10" & x"054" => data <= x"a0";
            when "10" & x"055" => data <= x"bd";
            when "10" & x"056" => data <= x"45";
            when "10" & x"057" => data <= x"0d";
            when "10" & x"058" => data <= x"20";
            when "10" & x"059" => data <= x"69";
            when "10" & x"05a" => data <= x"a0";
            when "10" & x"05b" => data <= x"bd";
            when "10" & x"05c" => data <= x"46";
            when "10" & x"05d" => data <= x"0d";
            when "10" & x"05e" => data <= x"20";
            when "10" & x"05f" => data <= x"69";
            when "10" & x"060" => data <= x"a0";
            when "10" & x"061" => data <= x"a9";
            when "10" & x"062" => data <= x"00";
            when "10" & x"063" => data <= x"99";
            when "10" & x"064" => data <= x"00";
            when "10" & x"065" => data <= x"01";
            when "10" & x"066" => data <= x"4c";
            when "10" & x"067" => data <= x"00";
            when "10" & x"068" => data <= x"01";
            when "10" & x"069" => data <= x"48";
            when "10" & x"06a" => data <= x"4a";
            when "10" & x"06b" => data <= x"4a";
            when "10" & x"06c" => data <= x"4a";
            when "10" & x"06d" => data <= x"4a";
            when "10" & x"06e" => data <= x"20";
            when "10" & x"06f" => data <= x"74";
            when "10" & x"070" => data <= x"a0";
            when "10" & x"071" => data <= x"68";
            when "10" & x"072" => data <= x"29";
            when "10" & x"073" => data <= x"0f";
            when "10" & x"074" => data <= x"18";
            when "10" & x"075" => data <= x"69";
            when "10" & x"076" => data <= x"30";
            when "10" & x"077" => data <= x"c9";
            when "10" & x"078" => data <= x"3a";
            when "10" & x"079" => data <= x"90";
            when "10" & x"07a" => data <= x"02";
            when "10" & x"07b" => data <= x"69";
            when "10" & x"07c" => data <= x"06";
            when "10" & x"07d" => data <= x"99";
            when "10" & x"07e" => data <= x"00";
            when "10" & x"07f" => data <= x"01";
            when "10" & x"080" => data <= x"c8";
            when "10" & x"081" => data <= x"60";
            when "10" & x"082" => data <= x"20";
            when "10" & x"083" => data <= x"00";
            when "10" & x"084" => data <= x"a0";
            when "10" & x"085" => data <= x"11";
            when "10" & x"086" => data <= x"45";
            when "10" & x"087" => data <= x"73";
            when "10" & x"088" => data <= x"63";
            when "10" & x"089" => data <= x"61";
            when "10" & x"08a" => data <= x"70";
            when "10" & x"08b" => data <= x"65";
            when "10" & x"08c" => data <= x"00";
            when "10" & x"08d" => data <= x"48";
            when "10" & x"08e" => data <= x"a9";
            when "10" & x"08f" => data <= x"ff";
            when "10" & x"090" => data <= x"8d";
            when "10" & x"091" => data <= x"74";
            when "10" & x"092" => data <= x"10";
            when "10" & x"093" => data <= x"8d";
            when "10" & x"094" => data <= x"75";
            when "10" & x"095" => data <= x"10";
            when "10" & x"096" => data <= x"68";
            when "10" & x"097" => data <= x"60";
            when "10" & x"098" => data <= x"48";
            when "10" & x"099" => data <= x"a5";
            when "10" & x"09a" => data <= x"be";
            when "10" & x"09b" => data <= x"8d";
            when "10" & x"09c" => data <= x"72";
            when "10" & x"09d" => data <= x"10";
            when "10" & x"09e" => data <= x"a5";
            when "10" & x"09f" => data <= x"bf";
            when "10" & x"0a0" => data <= x"8d";
            when "10" & x"0a1" => data <= x"73";
            when "10" & x"0a2" => data <= x"10";
            when "10" & x"0a3" => data <= x"ad";
            when "10" & x"0a4" => data <= x"74";
            when "10" & x"0a5" => data <= x"10";
            when "10" & x"0a6" => data <= x"2d";
            when "10" & x"0a7" => data <= x"75";
            when "10" & x"0a8" => data <= x"10";
            when "10" & x"0a9" => data <= x"0d";
            when "10" & x"0aa" => data <= x"d7";
            when "10" & x"0ab" => data <= x"10";
            when "10" & x"0ac" => data <= x"49";
            when "10" & x"0ad" => data <= x"ff";
            when "10" & x"0ae" => data <= x"8d";
            when "10" & x"0af" => data <= x"d6";
            when "10" & x"0b0" => data <= x"10";
            when "10" & x"0b1" => data <= x"38";
            when "10" & x"0b2" => data <= x"f0";
            when "10" & x"0b3" => data <= x"0d";
            when "10" & x"0b4" => data <= x"20";
            when "10" & x"0b5" => data <= x"c3";
            when "10" & x"0b6" => data <= x"a0";
            when "10" & x"0b7" => data <= x"a2";
            when "10" & x"0b8" => data <= x"72";
            when "10" & x"0b9" => data <= x"a0";
            when "10" & x"0ba" => data <= x"10";
            when "10" & x"0bb" => data <= x"68";
            when "10" & x"0bc" => data <= x"48";
            when "10" & x"0bd" => data <= x"20";
            when "10" & x"0be" => data <= x"06";
            when "10" & x"0bf" => data <= x"04";
            when "10" & x"0c0" => data <= x"18";
            when "10" & x"0c1" => data <= x"68";
            when "10" & x"0c2" => data <= x"60";
            when "10" & x"0c3" => data <= x"48";
            when "10" & x"0c4" => data <= x"a9";
            when "10" & x"0c5" => data <= x"c1";
            when "10" & x"0c6" => data <= x"20";
            when "10" & x"0c7" => data <= x"06";
            when "10" & x"0c8" => data <= x"04";
            when "10" & x"0c9" => data <= x"90";
            when "10" & x"0ca" => data <= x"f9";
            when "10" & x"0cb" => data <= x"68";
            when "10" & x"0cc" => data <= x"60";
            when "10" & x"0cd" => data <= x"ad";
            when "10" & x"0ce" => data <= x"d6";
            when "10" & x"0cf" => data <= x"10";
            when "10" & x"0d0" => data <= x"f0";
            when "10" & x"0d1" => data <= x"05";
            when "10" & x"0d2" => data <= x"a9";
            when "10" & x"0d3" => data <= x"81";
            when "10" & x"0d4" => data <= x"20";
            when "10" & x"0d5" => data <= x"06";
            when "10" & x"0d6" => data <= x"04";
            when "10" & x"0d7" => data <= x"60";
            when "10" & x"0d8" => data <= x"9d";
            when "10" & x"0d9" => data <= x"05";
            when "10" & x"0da" => data <= x"01";
            when "10" & x"0db" => data <= x"20";
            when "10" & x"0dc" => data <= x"e4";
            when "10" & x"0dd" => data <= x"95";
            when "10" & x"0de" => data <= x"08";
            when "10" & x"0df" => data <= x"ad";
            when "10" & x"0e0" => data <= x"81";
            when "10" & x"0e1" => data <= x"10";
            when "10" & x"0e2" => data <= x"f0";
            when "10" & x"0e3" => data <= x"05";
            when "10" & x"0e4" => data <= x"a9";
            when "10" & x"0e5" => data <= x"81";
            when "10" & x"0e6" => data <= x"20";
            when "10" & x"0e7" => data <= x"06";
            when "10" & x"0e8" => data <= x"04";
            when "10" & x"0e9" => data <= x"28";
            when "10" & x"0ea" => data <= x"60";
            when "10" & x"0eb" => data <= x"f0";
            when "10" & x"0ec" => data <= x"06";
            when "10" & x"0ed" => data <= x"20";
            when "10" & x"0ee" => data <= x"c3";
            when "10" & x"0ef" => data <= x"a0";
            when "10" & x"0f0" => data <= x"18";
            when "10" & x"0f1" => data <= x"a9";
            when "10" & x"0f2" => data <= x"ff";
            when "10" & x"0f3" => data <= x"4c";
            when "10" & x"0f4" => data <= x"17";
            when "10" & x"0f5" => data <= x"96";
            when "10" & x"0f6" => data <= x"c9";
            when "10" & x"0f7" => data <= x"fe";
            when "10" & x"0f8" => data <= x"90";
            when "10" & x"0f9" => data <= x"5a";
            when "10" & x"0fa" => data <= x"d0";
            when "10" & x"0fb" => data <= x"1b";
            when "10" & x"0fc" => data <= x"c0";
            when "10" & x"0fd" => data <= x"00";
            when "10" & x"0fe" => data <= x"f0";
            when "10" & x"0ff" => data <= x"54";
            when "10" & x"100" => data <= x"a2";
            when "10" & x"101" => data <= x"06";
            when "10" & x"102" => data <= x"a9";
            when "10" & x"103" => data <= x"14";
            when "10" & x"104" => data <= x"20";
            when "10" & x"105" => data <= x"f4";
            when "10" & x"106" => data <= x"ff";
            when "10" & x"107" => data <= x"2c";
            when "10" & x"108" => data <= x"e0";
            when "10" & x"109" => data <= x"fe";
            when "10" & x"10a" => data <= x"10";
            when "10" & x"10b" => data <= x"fb";
            when "10" & x"10c" => data <= x"ad";
            when "10" & x"10d" => data <= x"e1";
            when "10" & x"10e" => data <= x"fe";
            when "10" & x"10f" => data <= x"f0";
            when "10" & x"110" => data <= x"41";
            when "10" & x"111" => data <= x"20";
            when "10" & x"112" => data <= x"ee";
            when "10" & x"113" => data <= x"ff";
            when "10" & x"114" => data <= x"4c";
            when "10" & x"115" => data <= x"07";
            when "10" & x"116" => data <= x"a1";
            when "10" & x"117" => data <= x"a9";
            when "10" & x"118" => data <= x"ad";
            when "10" & x"119" => data <= x"8d";
            when "10" & x"11a" => data <= x"20";
            when "10" & x"11b" => data <= x"02";
            when "10" & x"11c" => data <= x"a9";
            when "10" & x"11d" => data <= x"06";
            when "10" & x"11e" => data <= x"8d";
            when "10" & x"11f" => data <= x"21";
            when "10" & x"120" => data <= x"02";
            when "10" & x"121" => data <= x"a9";
            when "10" & x"122" => data <= x"16";
            when "10" & x"123" => data <= x"8d";
            when "10" & x"124" => data <= x"02";
            when "10" & x"125" => data <= x"02";
            when "10" & x"126" => data <= x"a0";
            when "10" & x"127" => data <= x"00";
            when "10" & x"128" => data <= x"8c";
            when "10" & x"129" => data <= x"03";
            when "10" & x"12a" => data <= x"02";
            when "10" & x"12b" => data <= x"a9";
            when "10" & x"12c" => data <= x"8e";
            when "10" & x"12d" => data <= x"8d";
            when "10" & x"12e" => data <= x"e0";
            when "10" & x"12f" => data <= x"fe";
            when "10" & x"130" => data <= x"b9";
            when "10" & x"131" => data <= x"03";
            when "10" & x"132" => data <= x"8b";
            when "10" & x"133" => data <= x"99";
            when "10" & x"134" => data <= x"00";
            when "10" & x"135" => data <= x"04";
            when "10" & x"136" => data <= x"b9";
            when "10" & x"137" => data <= x"03";
            when "10" & x"138" => data <= x"8c";
            when "10" & x"139" => data <= x"99";
            when "10" & x"13a" => data <= x"00";
            when "10" & x"13b" => data <= x"05";
            when "10" & x"13c" => data <= x"b9";
            when "10" & x"13d" => data <= x"03";
            when "10" & x"13e" => data <= x"8d";
            when "10" & x"13f" => data <= x"99";
            when "10" & x"140" => data <= x"00";
            when "10" & x"141" => data <= x"06";
            when "10" & x"142" => data <= x"88";
            when "10" & x"143" => data <= x"d0";
            when "10" & x"144" => data <= x"eb";
            when "10" & x"145" => data <= x"20";
            when "10" & x"146" => data <= x"21";
            when "10" & x"147" => data <= x"04";
            when "10" & x"148" => data <= x"a2";
            when "10" & x"149" => data <= x"40";
            when "10" & x"14a" => data <= x"bd";
            when "10" & x"14b" => data <= x"c2";
            when "10" & x"14c" => data <= x"8a";
            when "10" & x"14d" => data <= x"95";
            when "10" & x"14e" => data <= x"16";
            when "10" & x"14f" => data <= x"ca";
            when "10" & x"150" => data <= x"10";
            when "10" & x"151" => data <= x"f8";
            when "10" & x"152" => data <= x"a9";
            when "10" & x"153" => data <= x"00";
            when "10" & x"154" => data <= x"60";
            when "10" & x"155" => data <= x"a9";
            when "10" & x"156" => data <= x"00";
            when "10" & x"157" => data <= x"8d";
            when "10" & x"158" => data <= x"04";
            when "10" & x"159" => data <= x"0d";
            when "10" & x"15a" => data <= x"a9";
            when "10" & x"15b" => data <= x"ff";
            when "10" & x"15c" => data <= x"8d";
            when "10" & x"15d" => data <= x"52";
            when "10" & x"15e" => data <= x"0d";
            when "10" & x"15f" => data <= x"48";
            when "10" & x"160" => data <= x"4c";
            when "10" & x"161" => data <= x"3b";
            when "10" & x"162" => data <= x"93";
            when "10" & x"163" => data <= x"b9";
            when "10" & x"164" => data <= x"14";
            when "10" & x"165" => data <= x"11";
            when "10" & x"166" => data <= x"99";
            when "10" & x"167" => data <= x"10";
            when "10" & x"168" => data <= x"11";
            when "10" & x"169" => data <= x"b9";
            when "10" & x"16a" => data <= x"15";
            when "10" & x"16b" => data <= x"11";
            when "10" & x"16c" => data <= x"99";
            when "10" & x"16d" => data <= x"11";
            when "10" & x"16e" => data <= x"11";
            when "10" & x"16f" => data <= x"b9";
            when "10" & x"170" => data <= x"16";
            when "10" & x"171" => data <= x"11";
            when "10" & x"172" => data <= x"99";
            when "10" & x"173" => data <= x"12";
            when "10" & x"174" => data <= x"11";
            when "10" & x"175" => data <= x"60";
            when "10" & x"176" => data <= x"60";
            when "10" & x"177" => data <= x"a2";
            when "10" & x"178" => data <= x"06";
            when "10" & x"179" => data <= x"8e";
            when "10" & x"17a" => data <= x"40";
            when "10" & x"17b" => data <= x"fe";
            when "10" & x"17c" => data <= x"e8";
            when "10" & x"17d" => data <= x"8e";
            when "10" & x"17e" => data <= x"40";
            when "10" & x"17f" => data <= x"fe";
            when "10" & x"180" => data <= x"60";
            when "10" & x"181" => data <= x"a9";
            when "10" & x"182" => data <= x"76";
            when "10" & x"183" => data <= x"ea";
            when "10" & x"184" => data <= x"ea";
            when "10" & x"185" => data <= x"ea";
            when "10" & x"186" => data <= x"ea";
            when "10" & x"187" => data <= x"ea";
            when "10" & x"188" => data <= x"ea";
            when "10" & x"189" => data <= x"60";
            when "10" & x"18a" => data <= x"48";
            when "10" & x"18b" => data <= x"68";
            when "10" & x"18c" => data <= x"20";
            when "10" & x"18d" => data <= x"85";
            when "10" & x"18e" => data <= x"a1";
            when "10" & x"18f" => data <= x"60";
            when "10" & x"190" => data <= x"ad";
            when "10" & x"191" => data <= x"bb";
            when "10" & x"192" => data <= x"fc";
            when "10" & x"193" => data <= x"8d";
            when "10" & x"194" => data <= x"3a";
            when "10" & x"195" => data <= x"0d";
            when "10" & x"196" => data <= x"ad";
            when "10" & x"197" => data <= x"b2";
            when "10" & x"198" => data <= x"fc";
            when "10" & x"199" => data <= x"8d";
            when "10" & x"19a" => data <= x"3b";
            when "10" & x"19b" => data <= x"0d";
            when "10" & x"19c" => data <= x"60";
            when "10" & x"19d" => data <= x"a9";
            when "10" & x"19e" => data <= x"08";
            when "10" & x"19f" => data <= x"8d";
            when "10" & x"1a0" => data <= x"bb";
            when "10" & x"1a1" => data <= x"fc";
            when "10" & x"1a2" => data <= x"ad";
            when "10" & x"1a3" => data <= x"b2";
            when "10" & x"1a4" => data <= x"fc";
            when "10" & x"1a5" => data <= x"4d";
            when "10" & x"1a6" => data <= x"4c";
            when "10" & x"1a7" => data <= x"0d";
            when "10" & x"1a8" => data <= x"0d";
            when "10" & x"1a9" => data <= x"4b";
            when "10" & x"1aa" => data <= x"0d";
            when "10" & x"1ab" => data <= x"8d";
            when "10" & x"1ac" => data <= x"b2";
            when "10" & x"1ad" => data <= x"fc";
            when "10" & x"1ae" => data <= x"ad";
            when "10" & x"1af" => data <= x"4b";
            when "10" & x"1b0" => data <= x"0d";
            when "10" & x"1b1" => data <= x"0d";
            when "10" & x"1b2" => data <= x"3f";
            when "10" & x"1b3" => data <= x"0d";
            when "10" & x"1b4" => data <= x"0d";
            when "10" & x"1b5" => data <= x"51";
            when "10" & x"1b6" => data <= x"0d";
            when "10" & x"1b7" => data <= x"8d";
            when "10" & x"1b8" => data <= x"b0";
            when "10" & x"1b9" => data <= x"fc";
            when "10" & x"1ba" => data <= x"ad";
            when "10" & x"1bb" => data <= x"ba";
            when "10" & x"1bc" => data <= x"fc";
            when "10" & x"1bd" => data <= x"60";
            when "10" & x"1be" => data <= x"ad";
            when "10" & x"1bf" => data <= x"bd";
            when "10" & x"1c0" => data <= x"fc";
            when "10" & x"1c1" => data <= x"29";
            when "10" & x"1c2" => data <= x"04";
            when "10" & x"1c3" => data <= x"f0";
            when "10" & x"1c4" => data <= x"f9";
            when "10" & x"1c5" => data <= x"60";
            when "10" & x"1c6" => data <= x"ad";
            when "10" & x"1c7" => data <= x"4c";
            when "10" & x"1c8" => data <= x"0d";
            when "10" & x"1c9" => data <= x"0d";
            when "10" & x"1ca" => data <= x"3f";
            when "10" & x"1cb" => data <= x"0d";
            when "10" & x"1cc" => data <= x"0d";
            when "10" & x"1cd" => data <= x"51";
            when "10" & x"1ce" => data <= x"0d";
            when "10" & x"1cf" => data <= x"8d";
            when "10" & x"1d0" => data <= x"b0";
            when "10" & x"1d1" => data <= x"fc";
            when "10" & x"1d2" => data <= x"ad";
            when "10" & x"1d3" => data <= x"3b";
            when "10" & x"1d4" => data <= x"0d";
            when "10" & x"1d5" => data <= x"8d";
            when "10" & x"1d6" => data <= x"b2";
            when "10" & x"1d7" => data <= x"fc";
            when "10" & x"1d8" => data <= x"ad";
            when "10" & x"1d9" => data <= x"3a";
            when "10" & x"1da" => data <= x"0d";
            when "10" & x"1db" => data <= x"8d";
            when "10" & x"1dc" => data <= x"bb";
            when "10" & x"1dd" => data <= x"fc";
            when "10" & x"1de" => data <= x"ad";
            when "10" & x"1df" => data <= x"ba";
            when "10" & x"1e0" => data <= x"fc";
            when "10" & x"1e1" => data <= x"60";
            when "10" & x"1e2" => data <= x"20";
            when "10" & x"1e3" => data <= x"90";
            when "10" & x"1e4" => data <= x"a1";
            when "10" & x"1e5" => data <= x"20";
            when "10" & x"1e6" => data <= x"9d";
            when "10" & x"1e7" => data <= x"a1";
            when "10" & x"1e8" => data <= x"20";
            when "10" & x"1e9" => data <= x"be";
            when "10" & x"1ea" => data <= x"a1";
            when "10" & x"1eb" => data <= x"20";
            when "10" & x"1ec" => data <= x"c6";
            when "10" & x"1ed" => data <= x"a1";
            when "10" & x"1ee" => data <= x"60";
            when "10" & x"1ef" => data <= x"20";
            when "10" & x"1f0" => data <= x"90";
            when "10" & x"1f1" => data <= x"a1";
            when "10" & x"1f2" => data <= x"20";
            when "10" & x"1f3" => data <= x"9d";
            when "10" & x"1f4" => data <= x"a1";
            when "10" & x"1f5" => data <= x"c0";
            when "10" & x"1f6" => data <= x"ff";
            when "10" & x"1f7" => data <= x"f0";
            when "10" & x"1f8" => data <= x"0b";
            when "10" & x"1f9" => data <= x"20";
            when "10" & x"1fa" => data <= x"be";
            when "10" & x"1fb" => data <= x"a1";
            when "10" & x"1fc" => data <= x"ad";
            when "10" & x"1fd" => data <= x"ba";
            when "10" & x"1fe" => data <= x"fc";
            when "10" & x"1ff" => data <= x"91";
            when "10" & x"200" => data <= x"a0";
            when "10" & x"201" => data <= x"c8";
            when "10" & x"202" => data <= x"d0";
            when "10" & x"203" => data <= x"f1";
            when "10" & x"204" => data <= x"20";
            when "10" & x"205" => data <= x"be";
            when "10" & x"206" => data <= x"a1";
            when "10" & x"207" => data <= x"20";
            when "10" & x"208" => data <= x"c6";
            when "10" & x"209" => data <= x"a1";
            when "10" & x"20a" => data <= x"91";
            when "10" & x"20b" => data <= x"a0";
            when "10" & x"20c" => data <= x"e8";
            when "10" & x"20d" => data <= x"c8";
            when "10" & x"20e" => data <= x"60";
            when "10" & x"20f" => data <= x"ad";
            when "10" & x"210" => data <= x"4b";
            when "10" & x"211" => data <= x"0d";
            when "10" & x"212" => data <= x"0d";
            when "10" & x"213" => data <= x"3f";
            when "10" & x"214" => data <= x"0d";
            when "10" & x"215" => data <= x"0d";
            when "10" & x"216" => data <= x"51";
            when "10" & x"217" => data <= x"0d";
            when "10" & x"218" => data <= x"aa";
            when "10" & x"219" => data <= x"ad";
            when "10" & x"21a" => data <= x"4c";
            when "10" & x"21b" => data <= x"0d";
            when "10" & x"21c" => data <= x"0d";
            when "10" & x"21d" => data <= x"3f";
            when "10" & x"21e" => data <= x"0d";
            when "10" & x"21f" => data <= x"0d";
            when "10" & x"220" => data <= x"51";
            when "10" & x"221" => data <= x"0d";
            when "10" & x"222" => data <= x"8e";
            when "10" & x"223" => data <= x"b0";
            when "10" & x"224" => data <= x"fc";
            when "10" & x"225" => data <= x"8d";
            when "10" & x"226" => data <= x"b0";
            when "10" & x"227" => data <= x"fc";
            when "10" & x"228" => data <= x"8e";
            when "10" & x"229" => data <= x"b0";
            when "10" & x"22a" => data <= x"fc";
            when "10" & x"22b" => data <= x"8d";
            when "10" & x"22c" => data <= x"b0";
            when "10" & x"22d" => data <= x"fc";
            when "10" & x"22e" => data <= x"8e";
            when "10" & x"22f" => data <= x"b0";
            when "10" & x"230" => data <= x"fc";
            when "10" & x"231" => data <= x"8d";
            when "10" & x"232" => data <= x"b0";
            when "10" & x"233" => data <= x"fc";
            when "10" & x"234" => data <= x"8e";
            when "10" & x"235" => data <= x"b0";
            when "10" & x"236" => data <= x"fc";
            when "10" & x"237" => data <= x"8d";
            when "10" & x"238" => data <= x"b0";
            when "10" & x"239" => data <= x"fc";
            when "10" & x"23a" => data <= x"8e";
            when "10" & x"23b" => data <= x"b0";
            when "10" & x"23c" => data <= x"fc";
            when "10" & x"23d" => data <= x"8d";
            when "10" & x"23e" => data <= x"b0";
            when "10" & x"23f" => data <= x"fc";
            when "10" & x"240" => data <= x"8e";
            when "10" & x"241" => data <= x"b0";
            when "10" & x"242" => data <= x"fc";
            when "10" & x"243" => data <= x"8d";
            when "10" & x"244" => data <= x"b0";
            when "10" & x"245" => data <= x"fc";
            when "10" & x"246" => data <= x"8e";
            when "10" & x"247" => data <= x"b0";
            when "10" & x"248" => data <= x"fc";
            when "10" & x"249" => data <= x"8d";
            when "10" & x"24a" => data <= x"b0";
            when "10" & x"24b" => data <= x"fc";
            when "10" & x"24c" => data <= x"8e";
            when "10" & x"24d" => data <= x"b0";
            when "10" & x"24e" => data <= x"fc";
            when "10" & x"24f" => data <= x"8d";
            when "10" & x"250" => data <= x"b0";
            when "10" & x"251" => data <= x"fc";
            when "10" & x"252" => data <= x"ad";
            when "10" & x"253" => data <= x"ba";
            when "10" & x"254" => data <= x"fc";
            when "10" & x"255" => data <= x"60";
            when "10" & x"256" => data <= x"a9";
            when "10" & x"257" => data <= x"18";
            when "10" & x"258" => data <= x"8d";
            when "10" & x"259" => data <= x"bb";
            when "10" & x"25a" => data <= x"fc";
            when "10" & x"25b" => data <= x"a9";
            when "10" & x"25c" => data <= x"1d";
            when "10" & x"25d" => data <= x"8d";
            when "10" & x"25e" => data <= x"b2";
            when "10" & x"25f" => data <= x"fc";
            when "10" & x"260" => data <= x"a9";
            when "10" & x"261" => data <= x"14";
            when "10" & x"262" => data <= x"8d";
            when "10" & x"263" => data <= x"b0";
            when "10" & x"264" => data <= x"fc";
            when "10" & x"265" => data <= x"60";
            when "10" & x"266" => data <= x"20";
            when "10" & x"267" => data <= x"90";
            when "10" & x"268" => data <= x"a1";
            when "10" & x"269" => data <= x"20";
            when "10" & x"26a" => data <= x"56";
            when "10" & x"26b" => data <= x"a2";
            when "10" & x"26c" => data <= x"68";
            when "10" & x"26d" => data <= x"8d";
            when "10" & x"26e" => data <= x"ba";
            when "10" & x"26f" => data <= x"fc";
            when "10" & x"270" => data <= x"20";
            when "10" & x"271" => data <= x"be";
            when "10" & x"272" => data <= x"a1";
            when "10" & x"273" => data <= x"20";
            when "10" & x"274" => data <= x"8a";
            when "10" & x"275" => data <= x"a1";
            when "10" & x"276" => data <= x"4c";
            when "10" & x"277" => data <= x"c6";
            when "10" & x"278" => data <= x"a1";
            when "10" & x"279" => data <= x"20";
            when "10" & x"27a" => data <= x"90";
            when "10" & x"27b" => data <= x"a1";
            when "10" & x"27c" => data <= x"20";
            when "10" & x"27d" => data <= x"56";
            when "10" & x"27e" => data <= x"a2";
            when "10" & x"27f" => data <= x"b1";
            when "10" & x"280" => data <= x"a0";
            when "10" & x"281" => data <= x"8d";
            when "10" & x"282" => data <= x"ba";
            when "10" & x"283" => data <= x"fc";
            when "10" & x"284" => data <= x"20";
            when "10" & x"285" => data <= x"be";
            when "10" & x"286" => data <= x"a1";
            when "10" & x"287" => data <= x"c8";
            when "10" & x"288" => data <= x"d0";
            when "10" & x"289" => data <= x"f5";
            when "10" & x"28a" => data <= x"4c";
            when "10" & x"28b" => data <= x"c6";
            when "10" & x"28c" => data <= x"a1";
            when "10" & x"28d" => data <= x"ad";
            when "10" & x"28e" => data <= x"3f";
            when "10" & x"28f" => data <= x"0d";
            when "10" & x"290" => data <= x"d0";
            when "10" & x"291" => data <= x"e7";
            when "10" & x"292" => data <= x"b1";
            when "10" & x"293" => data <= x"a0";
            when "10" & x"294" => data <= x"20";
            when "10" & x"295" => data <= x"9b";
            when "10" & x"296" => data <= x"a2";
            when "10" & x"297" => data <= x"c8";
            when "10" & x"298" => data <= x"d0";
            when "10" & x"299" => data <= x"f8";
            when "10" & x"29a" => data <= x"60";
            when "10" & x"29b" => data <= x"86";
            when "10" & x"29c" => data <= x"b0";
            when "10" & x"29d" => data <= x"ae";
            when "10" & x"29e" => data <= x"4a";
            when "10" & x"29f" => data <= x"0d";
            when "10" & x"2a0" => data <= x"18";
            when "10" & x"2a1" => data <= x"2a";
            when "10" & x"2a2" => data <= x"2a";
            when "10" & x"2a3" => data <= x"ca";
            when "10" & x"2a4" => data <= x"d0";
            when "10" & x"2a5" => data <= x"fb";
            when "10" & x"2a6" => data <= x"48";
            when "10" & x"2a7" => data <= x"2d";
            when "10" & x"2a8" => data <= x"4c";
            when "10" & x"2a9" => data <= x"0d";
            when "10" & x"2aa" => data <= x"0d";
            when "10" & x"2ab" => data <= x"3f";
            when "10" & x"2ac" => data <= x"0d";
            when "10" & x"2ad" => data <= x"0d";
            when "10" & x"2ae" => data <= x"51";
            when "10" & x"2af" => data <= x"0d";
            when "10" & x"2b0" => data <= x"8d";
            when "10" & x"2b1" => data <= x"b0";
            when "10" & x"2b2" => data <= x"fc";
            when "10" & x"2b3" => data <= x"0d";
            when "10" & x"2b4" => data <= x"4e";
            when "10" & x"2b5" => data <= x"0d";
            when "10" & x"2b6" => data <= x"8d";
            when "10" & x"2b7" => data <= x"b0";
            when "10" & x"2b8" => data <= x"fc";
            when "10" & x"2b9" => data <= x"68";
            when "10" & x"2ba" => data <= x"a2";
            when "10" & x"2bb" => data <= x"07";
            when "10" & x"2bc" => data <= x"2a";
            when "10" & x"2bd" => data <= x"48";
            when "10" & x"2be" => data <= x"2d";
            when "10" & x"2bf" => data <= x"4c";
            when "10" & x"2c0" => data <= x"0d";
            when "10" & x"2c1" => data <= x"0d";
            when "10" & x"2c2" => data <= x"3f";
            when "10" & x"2c3" => data <= x"0d";
            when "10" & x"2c4" => data <= x"0d";
            when "10" & x"2c5" => data <= x"51";
            when "10" & x"2c6" => data <= x"0d";
            when "10" & x"2c7" => data <= x"2d";
            when "10" & x"2c8" => data <= x"4d";
            when "10" & x"2c9" => data <= x"0d";
            when "10" & x"2ca" => data <= x"8d";
            when "10" & x"2cb" => data <= x"b0";
            when "10" & x"2cc" => data <= x"fc";
            when "10" & x"2cd" => data <= x"0d";
            when "10" & x"2ce" => data <= x"4e";
            when "10" & x"2cf" => data <= x"0d";
            when "10" & x"2d0" => data <= x"8d";
            when "10" & x"2d1" => data <= x"b0";
            when "10" & x"2d2" => data <= x"fc";
            when "10" & x"2d3" => data <= x"68";
            when "10" & x"2d4" => data <= x"ca";
            when "10" & x"2d5" => data <= x"d0";
            when "10" & x"2d6" => data <= x"e5";
            when "10" & x"2d7" => data <= x"a6";
            when "10" & x"2d8" => data <= x"b0";
            when "10" & x"2d9" => data <= x"60";
            when "10" & x"2da" => data <= x"2c";
            when "10" & x"2db" => data <= x"40";
            when "10" & x"2dc" => data <= x"0d";
            when "10" & x"2dd" => data <= x"30";
            when "10" & x"2de" => data <= x"47";
            when "10" & x"2df" => data <= x"ad";
            when "10" & x"2e0" => data <= x"4b";
            when "10" & x"2e1" => data <= x"0d";
            when "10" & x"2e2" => data <= x"0d";
            when "10" & x"2e3" => data <= x"3f";
            when "10" & x"2e4" => data <= x"0d";
            when "10" & x"2e5" => data <= x"0d";
            when "10" & x"2e6" => data <= x"51";
            when "10" & x"2e7" => data <= x"0d";
            when "10" & x"2e8" => data <= x"aa";
            when "10" & x"2e9" => data <= x"ad";
            when "10" & x"2ea" => data <= x"4c";
            when "10" & x"2eb" => data <= x"0d";
            when "10" & x"2ec" => data <= x"0d";
            when "10" & x"2ed" => data <= x"3f";
            when "10" & x"2ee" => data <= x"0d";
            when "10" & x"2ef" => data <= x"0d";
            when "10" & x"2f0" => data <= x"51";
            when "10" & x"2f1" => data <= x"0d";
            when "10" & x"2f2" => data <= x"8e";
            when "10" & x"2f3" => data <= x"b0";
            when "10" & x"2f4" => data <= x"fc";
            when "10" & x"2f5" => data <= x"8d";
            when "10" & x"2f6" => data <= x"b0";
            when "10" & x"2f7" => data <= x"fc";
            when "10" & x"2f8" => data <= x"8e";
            when "10" & x"2f9" => data <= x"b0";
            when "10" & x"2fa" => data <= x"fc";
            when "10" & x"2fb" => data <= x"8d";
            when "10" & x"2fc" => data <= x"b0";
            when "10" & x"2fd" => data <= x"fc";
            when "10" & x"2fe" => data <= x"8e";
            when "10" & x"2ff" => data <= x"b0";
            when "10" & x"300" => data <= x"fc";
            when "10" & x"301" => data <= x"8d";
            when "10" & x"302" => data <= x"b0";
            when "10" & x"303" => data <= x"fc";
            when "10" & x"304" => data <= x"8e";
            when "10" & x"305" => data <= x"b0";
            when "10" & x"306" => data <= x"fc";
            when "10" & x"307" => data <= x"8d";
            when "10" & x"308" => data <= x"b0";
            when "10" & x"309" => data <= x"fc";
            when "10" & x"30a" => data <= x"8e";
            when "10" & x"30b" => data <= x"b0";
            when "10" & x"30c" => data <= x"fc";
            when "10" & x"30d" => data <= x"8d";
            when "10" & x"30e" => data <= x"b0";
            when "10" & x"30f" => data <= x"fc";
            when "10" & x"310" => data <= x"8e";
            when "10" & x"311" => data <= x"b0";
            when "10" & x"312" => data <= x"fc";
            when "10" & x"313" => data <= x"8d";
            when "10" & x"314" => data <= x"b0";
            when "10" & x"315" => data <= x"fc";
            when "10" & x"316" => data <= x"8e";
            when "10" & x"317" => data <= x"b0";
            when "10" & x"318" => data <= x"fc";
            when "10" & x"319" => data <= x"8d";
            when "10" & x"31a" => data <= x"b0";
            when "10" & x"31b" => data <= x"fc";
            when "10" & x"31c" => data <= x"8e";
            when "10" & x"31d" => data <= x"b0";
            when "10" & x"31e" => data <= x"fc";
            when "10" & x"31f" => data <= x"8d";
            when "10" & x"320" => data <= x"b0";
            when "10" & x"321" => data <= x"fc";
            when "10" & x"322" => data <= x"88";
            when "10" & x"323" => data <= x"d0";
            when "10" & x"324" => data <= x"cd";
            when "10" & x"325" => data <= x"60";
            when "10" & x"326" => data <= x"a9";
            when "10" & x"327" => data <= x"ff";
            when "10" & x"328" => data <= x"8d";
            when "10" & x"329" => data <= x"28";
            when "10" & x"32a" => data <= x"fc";
            when "10" & x"32b" => data <= x"ea";
            when "10" & x"32c" => data <= x"ea";
            when "10" & x"32d" => data <= x"ea";
            when "10" & x"32e" => data <= x"88";
            when "10" & x"32f" => data <= x"d0";
            when "10" & x"330" => data <= x"f7";
            when "10" & x"331" => data <= x"60";
            when "10" & x"332" => data <= x"a2";
            when "10" & x"333" => data <= x"00";
            when "10" & x"334" => data <= x"2c";
            when "10" & x"335" => data <= x"40";
            when "10" & x"336" => data <= x"0d";
            when "10" & x"337" => data <= x"30";
            when "10" & x"338" => data <= x"46";
            when "10" & x"339" => data <= x"8e";
            when "10" & x"33a" => data <= x"41";
            when "10" & x"33b" => data <= x"0d";
            when "10" & x"33c" => data <= x"a0";
            when "10" & x"33d" => data <= x"07";
            when "10" & x"33e" => data <= x"bd";
            when "10" & x"33f" => data <= x"42";
            when "10" & x"340" => data <= x"0d";
            when "10" & x"341" => data <= x"20";
            when "10" & x"342" => data <= x"9b";
            when "10" & x"343" => data <= x"a2";
            when "10" & x"344" => data <= x"e8";
            when "10" & x"345" => data <= x"88";
            when "10" & x"346" => data <= x"d0";
            when "10" & x"347" => data <= x"f6";
            when "10" & x"348" => data <= x"20";
            when "10" & x"349" => data <= x"4e";
            when "10" & x"34a" => data <= x"a3";
            when "10" & x"34b" => data <= x"4c";
            when "10" & x"34c" => data <= x"28";
            when "10" & x"34d" => data <= x"a2";
            when "10" & x"34e" => data <= x"a0";
            when "10" & x"34f" => data <= x"00";
            when "10" & x"350" => data <= x"84";
            when "10" & x"351" => data <= x"b0";
            when "10" & x"352" => data <= x"ad";
            when "10" & x"353" => data <= x"4b";
            when "10" & x"354" => data <= x"0d";
            when "10" & x"355" => data <= x"0d";
            when "10" & x"356" => data <= x"3f";
            when "10" & x"357" => data <= x"0d";
            when "10" & x"358" => data <= x"0d";
            when "10" & x"359" => data <= x"51";
            when "10" & x"35a" => data <= x"0d";
            when "10" & x"35b" => data <= x"aa";
            when "10" & x"35c" => data <= x"ad";
            when "10" & x"35d" => data <= x"4c";
            when "10" & x"35e" => data <= x"0d";
            when "10" & x"35f" => data <= x"0d";
            when "10" & x"360" => data <= x"3f";
            when "10" & x"361" => data <= x"0d";
            when "10" & x"362" => data <= x"0d";
            when "10" & x"363" => data <= x"51";
            when "10" & x"364" => data <= x"0d";
            when "10" & x"365" => data <= x"a8";
            when "10" & x"366" => data <= x"c6";
            when "10" & x"367" => data <= x"b0";
            when "10" & x"368" => data <= x"f0";
            when "10" & x"369" => data <= x"0f";
            when "10" & x"36a" => data <= x"8e";
            when "10" & x"36b" => data <= x"b0";
            when "10" & x"36c" => data <= x"fc";
            when "10" & x"36d" => data <= x"8c";
            when "10" & x"36e" => data <= x"b0";
            when "10" & x"36f" => data <= x"fc";
            when "10" & x"370" => data <= x"ad";
            when "10" & x"371" => data <= x"ba";
            when "10" & x"372" => data <= x"fc";
            when "10" & x"373" => data <= x"29";
            when "10" & x"374" => data <= x"01";
            when "10" & x"375" => data <= x"d0";
            when "10" & x"376" => data <= x"ef";
            when "10" & x"377" => data <= x"98";
            when "10" & x"378" => data <= x"60";
            when "10" & x"379" => data <= x"ad";
            when "10" & x"37a" => data <= x"ba";
            when "10" & x"37b" => data <= x"fc";
            when "10" & x"37c" => data <= x"c9";
            when "10" & x"37d" => data <= x"00";
            when "10" & x"37e" => data <= x"60";
            when "10" & x"37f" => data <= x"8e";
            when "10" & x"380" => data <= x"41";
            when "10" & x"381" => data <= x"0d";
            when "10" & x"382" => data <= x"a0";
            when "10" & x"383" => data <= x"08";
            when "10" & x"384" => data <= x"bd";
            when "10" & x"385" => data <= x"42";
            when "10" & x"386" => data <= x"0d";
            when "10" & x"387" => data <= x"8d";
            when "10" & x"388" => data <= x"28";
            when "10" & x"389" => data <= x"fc";
            when "10" & x"38a" => data <= x"ea";
            when "10" & x"38b" => data <= x"ea";
            when "10" & x"38c" => data <= x"e8";
            when "10" & x"38d" => data <= x"88";
            when "10" & x"38e" => data <= x"d0";
            when "10" & x"38f" => data <= x"f4";
            when "10" & x"390" => data <= x"8d";
            when "10" & x"391" => data <= x"28";
            when "10" & x"392" => data <= x"fc";
            when "10" & x"393" => data <= x"20";
            when "10" & x"394" => data <= x"31";
            when "10" & x"395" => data <= x"a3";
            when "10" & x"396" => data <= x"ad";
            when "10" & x"397" => data <= x"28";
            when "10" & x"398" => data <= x"fc";
            when "10" & x"399" => data <= x"10";
            when "10" & x"39a" => data <= x"e3";
            when "10" & x"39b" => data <= x"88";
            when "10" & x"39c" => data <= x"d0";
            when "10" & x"39d" => data <= x"f5";
            when "10" & x"39e" => data <= x"4c";
            when "10" & x"39f" => data <= x"7c";
            when "10" & x"3a0" => data <= x"a3";
            when "10" & x"3a1" => data <= x"2c";
            when "10" & x"3a2" => data <= x"40";
            when "10" & x"3a3" => data <= x"0d";
            when "10" & x"3a4" => data <= x"30";
            when "10" & x"3a5" => data <= x"08";
            when "10" & x"3a6" => data <= x"20";
            when "10" & x"3a7" => data <= x"e2";
            when "10" & x"3a8" => data <= x"a1";
            when "10" & x"3a9" => data <= x"c9";
            when "10" & x"3aa" => data <= x"fe";
            when "10" & x"3ab" => data <= x"d0";
            when "10" & x"3ac" => data <= x"f9";
            when "10" & x"3ad" => data <= x"60";
            when "10" & x"3ae" => data <= x"a2";
            when "10" & x"3af" => data <= x"ff";
            when "10" & x"3b0" => data <= x"8e";
            when "10" & x"3b1" => data <= x"28";
            when "10" & x"3b2" => data <= x"fc";
            when "10" & x"3b3" => data <= x"20";
            when "10" & x"3b4" => data <= x"31";
            when "10" & x"3b5" => data <= x"a3";
            when "10" & x"3b6" => data <= x"ad";
            when "10" & x"3b7" => data <= x"28";
            when "10" & x"3b8" => data <= x"fc";
            when "10" & x"3b9" => data <= x"c9";
            when "10" & x"3ba" => data <= x"fe";
            when "10" & x"3bb" => data <= x"d0";
            when "10" & x"3bc" => data <= x"f3";
            when "10" & x"3bd" => data <= x"60";
            when "10" & x"3be" => data <= x"2c";
            when "10" & x"3bf" => data <= x"40";
            when "10" & x"3c0" => data <= x"0d";
            when "10" & x"3c1" => data <= x"30";
            when "10" & x"3c2" => data <= x"0d";
            when "10" & x"3c3" => data <= x"ac";
            when "10" & x"3c4" => data <= x"d6";
            when "10" & x"3c5" => data <= x"10";
            when "10" & x"3c6" => data <= x"d0";
            when "10" & x"3c7" => data <= x"03";
            when "10" & x"3c8" => data <= x"4c";
            when "10" & x"3c9" => data <= x"ef";
            when "10" & x"3ca" => data <= x"a1";
            when "10" & x"3cb" => data <= x"a0";
            when "10" & x"3cc" => data <= x"00";
            when "10" & x"3cd" => data <= x"4c";
            when "10" & x"3ce" => data <= x"0e";
            when "10" & x"3cf" => data <= x"a4";
            when "10" & x"3d0" => data <= x"a2";
            when "10" & x"3d1" => data <= x"ff";
            when "10" & x"3d2" => data <= x"8e";
            when "10" & x"3d3" => data <= x"28";
            when "10" & x"3d4" => data <= x"fc";
            when "10" & x"3d5" => data <= x"ac";
            when "10" & x"3d6" => data <= x"d6";
            when "10" & x"3d7" => data <= x"10";
            when "10" & x"3d8" => data <= x"d0";
            when "10" & x"3d9" => data <= x"16";
            when "10" & x"3da" => data <= x"ea";
            when "10" & x"3db" => data <= x"ea";
            when "10" & x"3dc" => data <= x"ea";
            when "10" & x"3dd" => data <= x"ad";
            when "10" & x"3de" => data <= x"28";
            when "10" & x"3df" => data <= x"fc";
            when "10" & x"3e0" => data <= x"8e";
            when "10" & x"3e1" => data <= x"28";
            when "10" & x"3e2" => data <= x"fc";
            when "10" & x"3e3" => data <= x"91";
            when "10" & x"3e4" => data <= x"a0";
            when "10" & x"3e5" => data <= x"c8";
            when "10" & x"3e6" => data <= x"c0";
            when "10" & x"3e7" => data <= x"ff";
            when "10" & x"3e8" => data <= x"d0";
            when "10" & x"3e9" => data <= x"f3";
            when "10" & x"3ea" => data <= x"ad";
            when "10" & x"3eb" => data <= x"28";
            when "10" & x"3ec" => data <= x"fc";
            when "10" & x"3ed" => data <= x"91";
            when "10" & x"3ee" => data <= x"a0";
            when "10" & x"3ef" => data <= x"60";
            when "10" & x"3f0" => data <= x"a0";
            when "10" & x"3f1" => data <= x"00";
            when "10" & x"3f2" => data <= x"4c";
            when "10" & x"3f3" => data <= x"3e";
            when "10" & x"3f4" => data <= x"a4";
            when "10" & x"3f5" => data <= x"2c";
            when "10" & x"3f6" => data <= x"40";
            when "10" & x"3f7" => data <= x"0d";
            when "10" & x"3f8" => data <= x"30";
            when "10" & x"3f9" => data <= x"1e";
            when "10" & x"3fa" => data <= x"ac";
            when "10" & x"3fb" => data <= x"d6";
            when "10" & x"3fc" => data <= x"10";
            when "10" & x"3fd" => data <= x"d0";
            when "10" & x"3fe" => data <= x"0c";
            when "10" & x"3ff" => data <= x"20";
            when "10" & x"400" => data <= x"e2";
            when "10" & x"401" => data <= x"a1";
            when "10" & x"402" => data <= x"91";
            when "10" & x"403" => data <= x"a0";
            when "10" & x"404" => data <= x"c8";
            when "10" & x"405" => data <= x"ce";
            when "10" & x"406" => data <= x"29";
            when "10" & x"407" => data <= x"0d";
            when "10" & x"408" => data <= x"d0";
            when "10" & x"409" => data <= x"f5";
            when "10" & x"40a" => data <= x"60";
            when "10" & x"40b" => data <= x"ac";
            when "10" & x"40c" => data <= x"29";
            when "10" & x"40d" => data <= x"0d";
            when "10" & x"40e" => data <= x"20";
            when "10" & x"40f" => data <= x"e2";
            when "10" & x"410" => data <= x"a1";
            when "10" & x"411" => data <= x"8d";
            when "10" & x"412" => data <= x"e5";
            when "10" & x"413" => data <= x"fe";
            when "10" & x"414" => data <= x"88";
            when "10" & x"415" => data <= x"d0";
            when "10" & x"416" => data <= x"f7";
            when "10" & x"417" => data <= x"60";
            when "10" & x"418" => data <= x"a2";
            when "10" & x"419" => data <= x"ff";
            when "10" & x"41a" => data <= x"8e";
            when "10" & x"41b" => data <= x"28";
            when "10" & x"41c" => data <= x"fc";
            when "10" & x"41d" => data <= x"ac";
            when "10" & x"41e" => data <= x"d6";
            when "10" & x"41f" => data <= x"10";
            when "10" & x"420" => data <= x"d0";
            when "10" & x"421" => data <= x"19";
            when "10" & x"422" => data <= x"ce";
            when "10" & x"423" => data <= x"29";
            when "10" & x"424" => data <= x"0d";
            when "10" & x"425" => data <= x"f0";
            when "10" & x"426" => data <= x"0e";
            when "10" & x"427" => data <= x"ad";
            when "10" & x"428" => data <= x"28";
            when "10" & x"429" => data <= x"fc";
            when "10" & x"42a" => data <= x"8e";
            when "10" & x"42b" => data <= x"28";
            when "10" & x"42c" => data <= x"fc";
            when "10" & x"42d" => data <= x"91";
            when "10" & x"42e" => data <= x"a0";
            when "10" & x"42f" => data <= x"c8";
            when "10" & x"430" => data <= x"ce";
            when "10" & x"431" => data <= x"29";
            when "10" & x"432" => data <= x"0d";
            when "10" & x"433" => data <= x"d0";
            when "10" & x"434" => data <= x"f2";
            when "10" & x"435" => data <= x"ad";
            when "10" & x"436" => data <= x"28";
            when "10" & x"437" => data <= x"fc";
            when "10" & x"438" => data <= x"91";
            when "10" & x"439" => data <= x"a0";
            when "10" & x"43a" => data <= x"60";
            when "10" & x"43b" => data <= x"ac";
            when "10" & x"43c" => data <= x"29";
            when "10" & x"43d" => data <= x"0d";
            when "10" & x"43e" => data <= x"88";
            when "10" & x"43f" => data <= x"f0";
            when "10" & x"440" => data <= x"1a";
            when "10" & x"441" => data <= x"ea";
            when "10" & x"442" => data <= x"ad";
            when "10" & x"443" => data <= x"28";
            when "10" & x"444" => data <= x"fc";
            when "10" & x"445" => data <= x"8e";
            when "10" & x"446" => data <= x"28";
            when "10" & x"447" => data <= x"fc";
            when "10" & x"448" => data <= x"8d";
            when "10" & x"449" => data <= x"e5";
            when "10" & x"44a" => data <= x"fe";
            when "10" & x"44b" => data <= x"20";
            when "10" & x"44c" => data <= x"31";
            when "10" & x"44d" => data <= x"a3";
            when "10" & x"44e" => data <= x"20";
            when "10" & x"44f" => data <= x"31";
            when "10" & x"450" => data <= x"a3";
            when "10" & x"451" => data <= x"ea";
            when "10" & x"452" => data <= x"ea";
            when "10" & x"453" => data <= x"ea";
            when "10" & x"454" => data <= x"88";
            when "10" & x"455" => data <= x"d0";
            when "10" & x"456" => data <= x"ea";
            when "10" & x"457" => data <= x"ea";
            when "10" & x"458" => data <= x"ea";
            when "10" & x"459" => data <= x"ea";
            when "10" & x"45a" => data <= x"ea";
            when "10" & x"45b" => data <= x"ad";
            when "10" & x"45c" => data <= x"28";
            when "10" & x"45d" => data <= x"fc";
            when "10" & x"45e" => data <= x"8d";
            when "10" & x"45f" => data <= x"e5";
            when "10" & x"460" => data <= x"fe";
            when "10" & x"461" => data <= x"60";
            when "10" & x"462" => data <= x"2c";
            when "10" & x"463" => data <= x"40";
            when "10" & x"464" => data <= x"0d";
            when "10" & x"465" => data <= x"30";
            when "10" & x"466" => data <= x"0c";
            when "10" & x"467" => data <= x"a0";
            when "10" & x"468" => data <= x"00";
            when "10" & x"469" => data <= x"20";
            when "10" & x"46a" => data <= x"e2";
            when "10" & x"46b" => data <= x"a1";
            when "10" & x"46c" => data <= x"99";
            when "10" & x"46d" => data <= x"00";
            when "10" & x"46e" => data <= x"0e";
            when "10" & x"46f" => data <= x"c8";
            when "10" & x"470" => data <= x"d0";
            when "10" & x"471" => data <= x"f7";
            when "10" & x"472" => data <= x"60";
            when "10" & x"473" => data <= x"a0";
            when "10" & x"474" => data <= x"00";
            when "10" & x"475" => data <= x"a2";
            when "10" & x"476" => data <= x"ff";
            when "10" & x"477" => data <= x"8e";
            when "10" & x"478" => data <= x"28";
            when "10" & x"479" => data <= x"fc";
            when "10" & x"47a" => data <= x"20";
            when "10" & x"47b" => data <= x"31";
            when "10" & x"47c" => data <= x"a3";
            when "10" & x"47d" => data <= x"ad";
            when "10" & x"47e" => data <= x"28";
            when "10" & x"47f" => data <= x"fc";
            when "10" & x"480" => data <= x"8e";
            when "10" & x"481" => data <= x"28";
            when "10" & x"482" => data <= x"fc";
            when "10" & x"483" => data <= x"99";
            when "10" & x"484" => data <= x"00";
            when "10" & x"485" => data <= x"0e";
            when "10" & x"486" => data <= x"c8";
            when "10" & x"487" => data <= x"c0";
            when "10" & x"488" => data <= x"ff";
            when "10" & x"489" => data <= x"d0";
            when "10" & x"48a" => data <= x"f2";
            when "10" & x"48b" => data <= x"ad";
            when "10" & x"48c" => data <= x"28";
            when "10" & x"48d" => data <= x"fc";
            when "10" & x"48e" => data <= x"99";
            when "10" & x"48f" => data <= x"00";
            when "10" & x"490" => data <= x"0e";
            when "10" & x"491" => data <= x"60";
            when "10" & x"492" => data <= x"2c";
            when "10" & x"493" => data <= x"40";
            when "10" & x"494" => data <= x"0d";
            when "10" & x"495" => data <= x"30";
            when "10" & x"496" => data <= x"0a";
            when "10" & x"497" => data <= x"a0";
            when "10" & x"498" => data <= x"02";
            when "10" & x"499" => data <= x"20";
            when "10" & x"49a" => data <= x"df";
            when "10" & x"49b" => data <= x"a2";
            when "10" & x"49c" => data <= x"a9";
            when "10" & x"49d" => data <= x"fe";
            when "10" & x"49e" => data <= x"4c";
            when "10" & x"49f" => data <= x"9b";
            when "10" & x"4a0" => data <= x"a2";
            when "10" & x"4a1" => data <= x"a2";
            when "10" & x"4a2" => data <= x"ff";
            when "10" & x"4a3" => data <= x"8e";
            when "10" & x"4a4" => data <= x"28";
            when "10" & x"4a5" => data <= x"fc";
            when "10" & x"4a6" => data <= x"20";
            when "10" & x"4a7" => data <= x"31";
            when "10" & x"4a8" => data <= x"a3";
            when "10" & x"4a9" => data <= x"8e";
            when "10" & x"4aa" => data <= x"28";
            when "10" & x"4ab" => data <= x"fc";
            when "10" & x"4ac" => data <= x"20";
            when "10" & x"4ad" => data <= x"31";
            when "10" & x"4ae" => data <= x"a3";
            when "10" & x"4af" => data <= x"ca";
            when "10" & x"4b0" => data <= x"8e";
            when "10" & x"4b1" => data <= x"28";
            when "10" & x"4b2" => data <= x"fc";
            when "10" & x"4b3" => data <= x"60";
            when "10" & x"4b4" => data <= x"a0";
            when "10" & x"4b5" => data <= x"02";
            when "10" & x"4b6" => data <= x"2c";
            when "10" & x"4b7" => data <= x"40";
            when "10" & x"4b8" => data <= x"0d";
            when "10" & x"4b9" => data <= x"30";
            when "10" & x"4ba" => data <= x"18";
            when "10" & x"4bb" => data <= x"20";
            when "10" & x"4bc" => data <= x"df";
            when "10" & x"4bd" => data <= x"a2";
            when "10" & x"4be" => data <= x"20";
            when "10" & x"4bf" => data <= x"4e";
            when "10" & x"4c0" => data <= x"a3";
            when "10" & x"4c1" => data <= x"20";
            when "10" & x"4c2" => data <= x"3a";
            when "10" & x"4c3" => data <= x"a2";
            when "10" & x"4c4" => data <= x"a8";
            when "10" & x"4c5" => data <= x"29";
            when "10" & x"4c6" => data <= x"1f";
            when "10" & x"4c7" => data <= x"c9";
            when "10" & x"4c8" => data <= x"05";
            when "10" & x"4c9" => data <= x"d0";
            when "10" & x"4ca" => data <= x"2b";
            when "10" & x"4cb" => data <= x"20";
            when "10" & x"4cc" => data <= x"e2";
            when "10" & x"4cd" => data <= x"a1";
            when "10" & x"4ce" => data <= x"c9";
            when "10" & x"4cf" => data <= x"ff";
            when "10" & x"4d0" => data <= x"d0";
            when "10" & x"4d1" => data <= x"f9";
            when "10" & x"4d2" => data <= x"60";
            when "10" & x"4d3" => data <= x"20";
            when "10" & x"4d4" => data <= x"26";
            when "10" & x"4d5" => data <= x"a3";
            when "10" & x"4d6" => data <= x"a2";
            when "10" & x"4d7" => data <= x"ff";
            when "10" & x"4d8" => data <= x"8e";
            when "10" & x"4d9" => data <= x"28";
            when "10" & x"4da" => data <= x"fc";
            when "10" & x"4db" => data <= x"20";
            when "10" & x"4dc" => data <= x"31";
            when "10" & x"4dd" => data <= x"a3";
            when "10" & x"4de" => data <= x"ad";
            when "10" & x"4df" => data <= x"28";
            when "10" & x"4e0" => data <= x"fc";
            when "10" & x"4e1" => data <= x"a8";
            when "10" & x"4e2" => data <= x"29";
            when "10" & x"4e3" => data <= x"1f";
            when "10" & x"4e4" => data <= x"c9";
            when "10" & x"4e5" => data <= x"05";
            when "10" & x"4e6" => data <= x"d0";
            when "10" & x"4e7" => data <= x"0e";
            when "10" & x"4e8" => data <= x"a9";
            when "10" & x"4e9" => data <= x"ff";
            when "10" & x"4ea" => data <= x"8e";
            when "10" & x"4eb" => data <= x"28";
            when "10" & x"4ec" => data <= x"fc";
            when "10" & x"4ed" => data <= x"20";
            when "10" & x"4ee" => data <= x"31";
            when "10" & x"4ef" => data <= x"a3";
            when "10" & x"4f0" => data <= x"cd";
            when "10" & x"4f1" => data <= x"28";
            when "10" & x"4f2" => data <= x"fc";
            when "10" & x"4f3" => data <= x"d0";
            when "10" & x"4f4" => data <= x"f5";
            when "10" & x"4f5" => data <= x"60";
            when "10" & x"4f6" => data <= x"98";
            when "10" & x"4f7" => data <= x"20";
            when "10" & x"4f8" => data <= x"1f";
            when "10" & x"4f9" => data <= x"a0";
            when "10" & x"4fa" => data <= x"c5";
            when "10" & x"4fb" => data <= x"4d";
            when "10" & x"4fc" => data <= x"4d";
            when "10" & x"4fd" => data <= x"43";
            when "10" & x"4fe" => data <= x"20";
            when "10" & x"4ff" => data <= x"57";
            when "10" & x"500" => data <= x"72";
            when "10" & x"501" => data <= x"69";
            when "10" & x"502" => data <= x"74";
            when "10" & x"503" => data <= x"65";
            when "10" & x"504" => data <= x"20";
            when "10" & x"505" => data <= x"72";
            when "10" & x"506" => data <= x"65";
            when "10" & x"507" => data <= x"73";
            when "10" & x"508" => data <= x"70";
            when "10" & x"509" => data <= x"6f";
            when "10" & x"50a" => data <= x"6e";
            when "10" & x"50b" => data <= x"73";
            when "10" & x"50c" => data <= x"65";
            when "10" & x"50d" => data <= x"20";
            when "10" & x"50e" => data <= x"66";
            when "10" & x"50f" => data <= x"61";
            when "10" & x"510" => data <= x"75";
            when "10" & x"511" => data <= x"6c";
            when "10" & x"512" => data <= x"74";
            when "10" & x"513" => data <= x"20";
            when "10" & x"514" => data <= x"00";
            when "10" & x"515" => data <= x"2c";
            when "10" & x"516" => data <= x"40";
            when "10" & x"517" => data <= x"0d";
            when "10" & x"518" => data <= x"30";
            when "10" & x"519" => data <= x"14";
            when "10" & x"51a" => data <= x"ac";
            when "10" & x"51b" => data <= x"d6";
            when "10" & x"51c" => data <= x"10";
            when "10" & x"51d" => data <= x"d0";
            when "10" & x"51e" => data <= x"03";
            when "10" & x"51f" => data <= x"4c";
            when "10" & x"520" => data <= x"8d";
            when "10" & x"521" => data <= x"a2";
            when "10" & x"522" => data <= x"a0";
            when "10" & x"523" => data <= x"00";
            when "10" & x"524" => data <= x"ad";
            when "10" & x"525" => data <= x"e5";
            when "10" & x"526" => data <= x"fe";
            when "10" & x"527" => data <= x"20";
            when "10" & x"528" => data <= x"9b";
            when "10" & x"529" => data <= x"a2";
            when "10" & x"52a" => data <= x"c8";
            when "10" & x"52b" => data <= x"d0";
            when "10" & x"52c" => data <= x"f7";
            when "10" & x"52d" => data <= x"60";
            when "10" & x"52e" => data <= x"ac";
            when "10" & x"52f" => data <= x"d6";
            when "10" & x"530" => data <= x"10";
            when "10" & x"531" => data <= x"d0";
            when "10" & x"532" => data <= x"09";
            when "10" & x"533" => data <= x"b1";
            when "10" & x"534" => data <= x"a0";
            when "10" & x"535" => data <= x"8d";
            when "10" & x"536" => data <= x"28";
            when "10" & x"537" => data <= x"fc";
            when "10" & x"538" => data <= x"c8";
            when "10" & x"539" => data <= x"d0";
            when "10" & x"53a" => data <= x"f8";
            when "10" & x"53b" => data <= x"60";
            when "10" & x"53c" => data <= x"a0";
            when "10" & x"53d" => data <= x"00";
            when "10" & x"53e" => data <= x"ad";
            when "10" & x"53f" => data <= x"e5";
            when "10" & x"540" => data <= x"fe";
            when "10" & x"541" => data <= x"8d";
            when "10" & x"542" => data <= x"28";
            when "10" & x"543" => data <= x"fc";
            when "10" & x"544" => data <= x"20";
            when "10" & x"545" => data <= x"31";
            when "10" & x"546" => data <= x"a3";
            when "10" & x"547" => data <= x"20";
            when "10" & x"548" => data <= x"31";
            when "10" & x"549" => data <= x"a3";
            when "10" & x"54a" => data <= x"20";
            when "10" & x"54b" => data <= x"31";
            when "10" & x"54c" => data <= x"a3";
            when "10" & x"54d" => data <= x"c8";
            when "10" & x"54e" => data <= x"d0";
            when "10" & x"54f" => data <= x"ee";
            when "10" & x"550" => data <= x"60";
            when "10" & x"551" => data <= x"2c";
            when "10" & x"552" => data <= x"40";
            when "10" & x"553" => data <= x"0d";
            when "10" & x"554" => data <= x"30";
            when "10" & x"555" => data <= x"0c";
            when "10" & x"556" => data <= x"a0";
            when "10" & x"557" => data <= x"00";
            when "10" & x"558" => data <= x"b9";
            when "10" & x"559" => data <= x"00";
            when "10" & x"55a" => data <= x"0e";
            when "10" & x"55b" => data <= x"20";
            when "10" & x"55c" => data <= x"9b";
            when "10" & x"55d" => data <= x"a2";
            when "10" & x"55e" => data <= x"c8";
            when "10" & x"55f" => data <= x"d0";
            when "10" & x"560" => data <= x"f7";
            when "10" & x"561" => data <= x"60";
            when "10" & x"562" => data <= x"a0";
            when "10" & x"563" => data <= x"00";
            when "10" & x"564" => data <= x"ea";
            when "10" & x"565" => data <= x"b9";
            when "10" & x"566" => data <= x"00";
            when "10" & x"567" => data <= x"0e";
            when "10" & x"568" => data <= x"8d";
            when "10" & x"569" => data <= x"28";
            when "10" & x"56a" => data <= x"fc";
            when "10" & x"56b" => data <= x"c8";
            when "10" & x"56c" => data <= x"d0";
            when "10" & x"56d" => data <= x"f6";
            when "10" & x"56e" => data <= x"60";
            when "10" & x"56f" => data <= x"a2";
            when "10" & x"570" => data <= x"00";
            when "10" & x"571" => data <= x"9d";
            when "10" & x"572" => data <= x"43";
            when "10" & x"573" => data <= x"0d";
            when "10" & x"574" => data <= x"a9";
            when "10" & x"575" => data <= x"00";
            when "10" & x"576" => data <= x"9d";
            when "10" & x"577" => data <= x"44";
            when "10" & x"578" => data <= x"0d";
            when "10" & x"579" => data <= x"9d";
            when "10" & x"57a" => data <= x"45";
            when "10" & x"57b" => data <= x"0d";
            when "10" & x"57c" => data <= x"9d";
            when "10" & x"57d" => data <= x"46";
            when "10" & x"57e" => data <= x"0d";
            when "10" & x"57f" => data <= x"9d";
            when "10" & x"580" => data <= x"47";
            when "10" & x"581" => data <= x"0d";
            when "10" & x"582" => data <= x"a9";
            when "10" & x"583" => data <= x"ff";
            when "10" & x"584" => data <= x"9d";
            when "10" & x"585" => data <= x"42";
            when "10" & x"586" => data <= x"0d";
            when "10" & x"587" => data <= x"9d";
            when "10" & x"588" => data <= x"48";
            when "10" & x"589" => data <= x"0d";
            when "10" & x"58a" => data <= x"9d";
            when "10" & x"58b" => data <= x"49";
            when "10" & x"58c" => data <= x"0d";
            when "10" & x"58d" => data <= x"ae";
            when "10" & x"58e" => data <= x"03";
            when "10" & x"58f" => data <= x"0d";
            when "10" & x"590" => data <= x"bd";
            when "10" & x"591" => data <= x"ae";
            when "10" & x"592" => data <= x"a5";
            when "10" & x"593" => data <= x"8d";
            when "10" & x"594" => data <= x"40";
            when "10" & x"595" => data <= x"0d";
            when "10" & x"596" => data <= x"60";
            when "10" & x"597" => data <= x"2c";
            when "10" & x"598" => data <= x"c9";
            when "10" & x"599" => data <= x"10";
            when "10" & x"59a" => data <= x"30";
            when "10" & x"59b" => data <= x"11";
            when "10" & x"59c" => data <= x"a9";
            when "10" & x"59d" => data <= x"8f";
            when "10" & x"59e" => data <= x"a2";
            when "10" & x"59f" => data <= x"0c";
            when "10" & x"5a0" => data <= x"a0";
            when "10" & x"5a1" => data <= x"ff";
            when "10" & x"5a2" => data <= x"20";
            when "10" & x"5a3" => data <= x"f4";
            when "10" & x"5a4" => data <= x"ff";
            when "10" & x"5a5" => data <= x"8c";
            when "10" & x"5a6" => data <= x"01";
            when "10" & x"5a7" => data <= x"0d";
            when "10" & x"5a8" => data <= x"a9";
            when "10" & x"5a9" => data <= x"ff";
            when "10" & x"5aa" => data <= x"8d";
            when "10" & x"5ab" => data <= x"c9";
            when "10" & x"5ac" => data <= x"10";
            when "10" & x"5ad" => data <= x"60";
            when "10" & x"5ae" => data <= x"00";
            when "10" & x"5af" => data <= x"80";
            when "10" & x"5b0" => data <= x"ad";
            when "10" & x"5b1" => data <= x"4f";
            when "10" & x"5b2" => data <= x"0d";
            when "10" & x"5b3" => data <= x"f0";
            when "10" & x"5b4" => data <= x"15";
            when "10" & x"5b5" => data <= x"ad";
            when "10" & x"5b6" => data <= x"3f";
            when "10" & x"5b7" => data <= x"0d";
            when "10" & x"5b8" => data <= x"d0";
            when "10" & x"5b9" => data <= x"26";
            when "10" & x"5ba" => data <= x"ad";
            when "10" & x"5bb" => data <= x"50";
            when "10" & x"5bc" => data <= x"0d";
            when "10" & x"5bd" => data <= x"d0";
            when "10" & x"5be" => data <= x"0b";
            when "10" & x"5bf" => data <= x"ad";
            when "10" & x"5c0" => data <= x"b2";
            when "10" & x"5c1" => data <= x"fc";
            when "10" & x"5c2" => data <= x"cd";
            when "10" & x"5c3" => data <= x"4c";
            when "10" & x"5c4" => data <= x"0d";
            when "10" & x"5c5" => data <= x"f0";
            when "10" & x"5c6" => data <= x"03";
            when "10" & x"5c7" => data <= x"20";
            when "10" & x"5c8" => data <= x"d6";
            when "10" & x"5c9" => data <= x"a9";
            when "10" & x"5ca" => data <= x"ad";
            when "10" & x"5cb" => data <= x"4c";
            when "10" & x"5cc" => data <= x"0d";
            when "10" & x"5cd" => data <= x"2d";
            when "10" & x"5ce" => data <= x"50";
            when "10" & x"5cf" => data <= x"0d";
            when "10" & x"5d0" => data <= x"d0";
            when "10" & x"5d1" => data <= x"36";
            when "10" & x"5d2" => data <= x"ad";
            when "10" & x"5d3" => data <= x"4c";
            when "10" & x"5d4" => data <= x"0d";
            when "10" & x"5d5" => data <= x"0d";
            when "10" & x"5d6" => data <= x"50";
            when "10" & x"5d7" => data <= x"0d";
            when "10" & x"5d8" => data <= x"8d";
            when "10" & x"5d9" => data <= x"b2";
            when "10" & x"5da" => data <= x"fc";
            when "10" & x"5db" => data <= x"ad";
            when "10" & x"5dc" => data <= x"3f";
            when "10" & x"5dd" => data <= x"0d";
            when "10" & x"5de" => data <= x"f0";
            when "10" & x"5df" => data <= x"0a";
            when "10" & x"5e0" => data <= x"a9";
            when "10" & x"5e1" => data <= x"1f";
            when "10" & x"5e2" => data <= x"8d";
            when "10" & x"5e3" => data <= x"b2";
            when "10" & x"5e4" => data <= x"fc";
            when "10" & x"5e5" => data <= x"a9";
            when "10" & x"5e6" => data <= x"00";
            when "10" & x"5e7" => data <= x"8d";
            when "10" & x"5e8" => data <= x"50";
            when "10" & x"5e9" => data <= x"0d";
            when "10" & x"5ea" => data <= x"ad";
            when "10" & x"5eb" => data <= x"3f";
            when "10" & x"5ec" => data <= x"0d";
            when "10" & x"5ed" => data <= x"d0";
            when "10" & x"5ee" => data <= x"03";
            when "10" & x"5ef" => data <= x"0d";
            when "10" & x"5f0" => data <= x"51";
            when "10" & x"5f1" => data <= x"0d";
            when "10" & x"5f2" => data <= x"8d";
            when "10" & x"5f3" => data <= x"b0";
            when "10" & x"5f4" => data <= x"fc";
            when "10" & x"5f5" => data <= x"ad";
            when "10" & x"5f6" => data <= x"bb";
            when "10" & x"5f7" => data <= x"fc";
            when "10" & x"5f8" => data <= x"29";
            when "10" & x"5f9" => data <= x"e3";
            when "10" & x"5fa" => data <= x"8d";
            when "10" & x"5fb" => data <= x"bb";
            when "10" & x"5fc" => data <= x"fc";
            when "10" & x"5fd" => data <= x"a9";
            when "10" & x"5fe" => data <= x"1c";
            when "10" & x"5ff" => data <= x"8d";
            when "10" & x"600" => data <= x"be";
            when "10" & x"601" => data <= x"fc";
            when "10" & x"602" => data <= x"a9";
            when "10" & x"603" => data <= x"00";
            when "10" & x"604" => data <= x"8d";
            when "10" & x"605" => data <= x"ba";
            when "10" & x"606" => data <= x"fc";
            when "10" & x"607" => data <= x"60";
            when "10" & x"608" => data <= x"20";
            when "10" & x"609" => data <= x"00";
            when "10" & x"60a" => data <= x"a0";
            when "10" & x"60b" => data <= x"ff";
            when "10" & x"60c" => data <= x"55";
            when "10" & x"60d" => data <= x"73";
            when "10" & x"60e" => data <= x"65";
            when "10" & x"60f" => data <= x"72";
            when "10" & x"610" => data <= x"20";
            when "10" & x"611" => data <= x"70";
            when "10" & x"612" => data <= x"6f";
            when "10" & x"613" => data <= x"72";
            when "10" & x"614" => data <= x"74";
            when "10" & x"615" => data <= x"20";
            when "10" & x"616" => data <= x"63";
            when "10" & x"617" => data <= x"6f";
            when "10" & x"618" => data <= x"6e";
            when "10" & x"619" => data <= x"66";
            when "10" & x"61a" => data <= x"6c";
            when "10" & x"61b" => data <= x"69";
            when "10" & x"61c" => data <= x"63";
            when "10" & x"61d" => data <= x"74";
            when "10" & x"61e" => data <= x"00";
            when "10" & x"61f" => data <= x"ad";
            when "10" & x"620" => data <= x"02";
            when "10" & x"621" => data <= x"0d";
            when "10" & x"622" => data <= x"c9";
            when "10" & x"623" => data <= x"54";
            when "10" & x"624" => data <= x"d0";
            when "10" & x"625" => data <= x"04";
            when "10" & x"626" => data <= x"20";
            when "10" & x"627" => data <= x"b0";
            when "10" & x"628" => data <= x"a5";
            when "10" & x"629" => data <= x"60";
            when "10" & x"62a" => data <= x"20";
            when "10" & x"62b" => data <= x"43";
            when "10" & x"62c" => data <= x"a6";
            when "10" & x"62d" => data <= x"d0";
            when "10" & x"62e" => data <= x"fa";
            when "10" & x"62f" => data <= x"20";
            when "10" & x"630" => data <= x"eb";
            when "10" & x"631" => data <= x"a9";
            when "10" & x"632" => data <= x"c9";
            when "10" & x"633" => data <= x"ff";
            when "10" & x"634" => data <= x"f0";
            when "10" & x"635" => data <= x"f3";
            when "10" & x"636" => data <= x"20";
            when "10" & x"637" => data <= x"00";
            when "10" & x"638" => data <= x"a0";
            when "10" & x"639" => data <= x"ff";
            when "10" & x"63a" => data <= x"43";
            when "10" & x"63b" => data <= x"61";
            when "10" & x"63c" => data <= x"72";
            when "10" & x"63d" => data <= x"64";
            when "10" & x"63e" => data <= x"3f";
            when "10" & x"63f" => data <= x"00";
            when "10" & x"640" => data <= x"20";
            when "10" & x"641" => data <= x"76";
            when "10" & x"642" => data <= x"a1";
            when "10" & x"643" => data <= x"20";
            when "10" & x"644" => data <= x"b0";
            when "10" & x"645" => data <= x"a5";
            when "10" & x"646" => data <= x"a0";
            when "10" & x"647" => data <= x"0a";
            when "10" & x"648" => data <= x"20";
            when "10" & x"649" => data <= x"da";
            when "10" & x"64a" => data <= x"a2";
            when "10" & x"64b" => data <= x"a9";
            when "10" & x"64c" => data <= x"40";
            when "10" & x"64d" => data <= x"20";
            when "10" & x"64e" => data <= x"6f";
            when "10" & x"64f" => data <= x"a5";
            when "10" & x"650" => data <= x"a9";
            when "10" & x"651" => data <= x"95";
            when "10" & x"652" => data <= x"8d";
            when "10" & x"653" => data <= x"48";
            when "10" & x"654" => data <= x"0d";
            when "10" & x"655" => data <= x"20";
            when "10" & x"656" => data <= x"32";
            when "10" & x"657" => data <= x"a3";
            when "10" & x"658" => data <= x"c9";
            when "10" & x"659" => data <= x"01";
            when "10" & x"65a" => data <= x"f0";
            when "10" & x"65b" => data <= x"03";
            when "10" & x"65c" => data <= x"4c";
            when "10" & x"65d" => data <= x"07";
            when "10" & x"65e" => data <= x"a7";
            when "10" & x"65f" => data <= x"a9";
            when "10" & x"660" => data <= x"01";
            when "10" & x"661" => data <= x"8d";
            when "10" & x"662" => data <= x"4f";
            when "10" & x"663" => data <= x"0d";
            when "10" & x"664" => data <= x"a9";
            when "10" & x"665" => data <= x"48";
            when "10" & x"666" => data <= x"20";
            when "10" & x"667" => data <= x"6f";
            when "10" & x"668" => data <= x"a5";
            when "10" & x"669" => data <= x"a9";
            when "10" & x"66a" => data <= x"01";
            when "10" & x"66b" => data <= x"8d";
            when "10" & x"66c" => data <= x"46";
            when "10" & x"66d" => data <= x"0d";
            when "10" & x"66e" => data <= x"a9";
            when "10" & x"66f" => data <= x"aa";
            when "10" & x"670" => data <= x"8d";
            when "10" & x"671" => data <= x"47";
            when "10" & x"672" => data <= x"0d";
            when "10" & x"673" => data <= x"a9";
            when "10" & x"674" => data <= x"87";
            when "10" & x"675" => data <= x"8d";
            when "10" & x"676" => data <= x"48";
            when "10" & x"677" => data <= x"0d";
            when "10" & x"678" => data <= x"20";
            when "10" & x"679" => data <= x"32";
            when "10" & x"67a" => data <= x"a3";
            when "10" & x"67b" => data <= x"c9";
            when "10" & x"67c" => data <= x"01";
            when "10" & x"67d" => data <= x"f0";
            when "10" & x"67e" => data <= x"20";
            when "10" & x"67f" => data <= x"a9";
            when "10" & x"680" => data <= x"02";
            when "10" & x"681" => data <= x"8d";
            when "10" & x"682" => data <= x"4f";
            when "10" & x"683" => data <= x"0d";
            when "10" & x"684" => data <= x"a9";
            when "10" & x"685" => data <= x"41";
            when "10" & x"686" => data <= x"20";
            when "10" & x"687" => data <= x"6f";
            when "10" & x"688" => data <= x"a5";
            when "10" & x"689" => data <= x"20";
            when "10" & x"68a" => data <= x"32";
            when "10" & x"68b" => data <= x"a3";
            when "10" & x"68c" => data <= x"c9";
            when "10" & x"68d" => data <= x"02";
            when "10" & x"68e" => data <= x"90";
            when "10" & x"68f" => data <= x"03";
            when "10" & x"690" => data <= x"4c";
            when "10" & x"691" => data <= x"07";
            when "10" & x"692" => data <= x"a7";
            when "10" & x"693" => data <= x"c9";
            when "10" & x"694" => data <= x"00";
            when "10" & x"695" => data <= x"d0";
            when "10" & x"696" => data <= x"ed";
            when "10" & x"697" => data <= x"a9";
            when "10" & x"698" => data <= x"02";
            when "10" & x"699" => data <= x"8d";
            when "10" & x"69a" => data <= x"4f";
            when "10" & x"69b" => data <= x"0d";
            when "10" & x"69c" => data <= x"4c";
            when "10" & x"69d" => data <= x"e7";
            when "10" & x"69e" => data <= x"a6";
            when "10" & x"69f" => data <= x"20";
            when "10" & x"6a0" => data <= x"e2";
            when "10" & x"6a1" => data <= x"a1";
            when "10" & x"6a2" => data <= x"20";
            when "10" & x"6a3" => data <= x"e2";
            when "10" & x"6a4" => data <= x"a1";
            when "10" & x"6a5" => data <= x"20";
            when "10" & x"6a6" => data <= x"e2";
            when "10" & x"6a7" => data <= x"a1";
            when "10" & x"6a8" => data <= x"20";
            when "10" & x"6a9" => data <= x"e2";
            when "10" & x"6aa" => data <= x"a1";
            when "10" & x"6ab" => data <= x"a9";
            when "10" & x"6ac" => data <= x"77";
            when "10" & x"6ad" => data <= x"20";
            when "10" & x"6ae" => data <= x"6f";
            when "10" & x"6af" => data <= x"a5";
            when "10" & x"6b0" => data <= x"20";
            when "10" & x"6b1" => data <= x"32";
            when "10" & x"6b2" => data <= x"a3";
            when "10" & x"6b3" => data <= x"a9";
            when "10" & x"6b4" => data <= x"69";
            when "10" & x"6b5" => data <= x"20";
            when "10" & x"6b6" => data <= x"6f";
            when "10" & x"6b7" => data <= x"a5";
            when "10" & x"6b8" => data <= x"a9";
            when "10" & x"6b9" => data <= x"40";
            when "10" & x"6ba" => data <= x"8d";
            when "10" & x"6bb" => data <= x"44";
            when "10" & x"6bc" => data <= x"0d";
            when "10" & x"6bd" => data <= x"20";
            when "10" & x"6be" => data <= x"32";
            when "10" & x"6bf" => data <= x"a3";
            when "10" & x"6c0" => data <= x"c9";
            when "10" & x"6c1" => data <= x"00";
            when "10" & x"6c2" => data <= x"d0";
            when "10" & x"6c3" => data <= x"e7";
            when "10" & x"6c4" => data <= x"a9";
            when "10" & x"6c5" => data <= x"7a";
            when "10" & x"6c6" => data <= x"20";
            when "10" & x"6c7" => data <= x"6f";
            when "10" & x"6c8" => data <= x"a5";
            when "10" & x"6c9" => data <= x"20";
            when "10" & x"6ca" => data <= x"32";
            when "10" & x"6cb" => data <= x"a3";
            when "10" & x"6cc" => data <= x"c9";
            when "10" & x"6cd" => data <= x"00";
            when "10" & x"6ce" => data <= x"d0";
            when "10" & x"6cf" => data <= x"37";
            when "10" & x"6d0" => data <= x"20";
            when "10" & x"6d1" => data <= x"e2";
            when "10" & x"6d2" => data <= x"a1";
            when "10" & x"6d3" => data <= x"29";
            when "10" & x"6d4" => data <= x"40";
            when "10" & x"6d5" => data <= x"48";
            when "10" & x"6d6" => data <= x"20";
            when "10" & x"6d7" => data <= x"e2";
            when "10" & x"6d8" => data <= x"a1";
            when "10" & x"6d9" => data <= x"20";
            when "10" & x"6da" => data <= x"e2";
            when "10" & x"6db" => data <= x"a1";
            when "10" & x"6dc" => data <= x"20";
            when "10" & x"6dd" => data <= x"e2";
            when "10" & x"6de" => data <= x"a1";
            when "10" & x"6df" => data <= x"68";
            when "10" & x"6e0" => data <= x"d0";
            when "10" & x"6e1" => data <= x"05";
            when "10" & x"6e2" => data <= x"a9";
            when "10" & x"6e3" => data <= x"02";
            when "10" & x"6e4" => data <= x"8d";
            when "10" & x"6e5" => data <= x"4f";
            when "10" & x"6e6" => data <= x"0d";
            when "10" & x"6e7" => data <= x"a9";
            when "10" & x"6e8" => data <= x"50";
            when "10" & x"6e9" => data <= x"20";
            when "10" & x"6ea" => data <= x"6f";
            when "10" & x"6eb" => data <= x"a5";
            when "10" & x"6ec" => data <= x"a9";
            when "10" & x"6ed" => data <= x"02";
            when "10" & x"6ee" => data <= x"8d";
            when "10" & x"6ef" => data <= x"46";
            when "10" & x"6f0" => data <= x"0d";
            when "10" & x"6f1" => data <= x"20";
            when "10" & x"6f2" => data <= x"32";
            when "10" & x"6f3" => data <= x"a3";
            when "10" & x"6f4" => data <= x"d0";
            when "10" & x"6f5" => data <= x"2e";
            when "10" & x"6f6" => data <= x"a9";
            when "10" & x"6f7" => data <= x"54";
            when "10" & x"6f8" => data <= x"8d";
            when "10" & x"6f9" => data <= x"02";
            when "10" & x"6fa" => data <= x"0d";
            when "10" & x"6fb" => data <= x"ad";
            when "10" & x"6fc" => data <= x"03";
            when "10" & x"6fd" => data <= x"0d";
            when "10" & x"6fe" => data <= x"8d";
            when "10" & x"6ff" => data <= x"04";
            when "10" & x"700" => data <= x"0d";
            when "10" & x"701" => data <= x"20";
            when "10" & x"702" => data <= x"80";
            when "10" & x"703" => data <= x"a1";
            when "10" & x"704" => data <= x"a9";
            when "10" & x"705" => data <= x"ff";
            when "10" & x"706" => data <= x"60";
            when "10" & x"707" => data <= x"ae";
            when "10" & x"708" => data <= x"03";
            when "10" & x"709" => data <= x"0d";
            when "10" & x"70a" => data <= x"e8";
            when "10" & x"70b" => data <= x"e0";
            when "10" & x"70c" => data <= x"02";
            when "10" & x"70d" => data <= x"b0";
            when "10" & x"70e" => data <= x"09";
            when "10" & x"70f" => data <= x"8e";
            when "10" & x"710" => data <= x"03";
            when "10" & x"711" => data <= x"0d";
            when "10" & x"712" => data <= x"20";
            when "10" & x"713" => data <= x"8d";
            when "10" & x"714" => data <= x"a5";
            when "10" & x"715" => data <= x"4c";
            when "10" & x"716" => data <= x"46";
            when "10" & x"717" => data <= x"a6";
            when "10" & x"718" => data <= x"a9";
            when "10" & x"719" => data <= x"00";
            when "10" & x"71a" => data <= x"8d";
            when "10" & x"71b" => data <= x"03";
            when "10" & x"71c" => data <= x"0d";
            when "10" & x"71d" => data <= x"20";
            when "10" & x"71e" => data <= x"8d";
            when "10" & x"71f" => data <= x"a5";
            when "10" & x"720" => data <= x"8d";
            when "10" & x"721" => data <= x"02";
            when "10" & x"722" => data <= x"0d";
            when "10" & x"723" => data <= x"60";
            when "10" & x"724" => data <= x"20";
            when "10" & x"725" => data <= x"1f";
            when "10" & x"726" => data <= x"a0";
            when "10" & x"727" => data <= x"ff";
            when "10" & x"728" => data <= x"53";
            when "10" & x"729" => data <= x"65";
            when "10" & x"72a" => data <= x"74";
            when "10" & x"72b" => data <= x"20";
            when "10" & x"72c" => data <= x"62";
            when "10" & x"72d" => data <= x"6c";
            when "10" & x"72e" => data <= x"6f";
            when "10" & x"72f" => data <= x"63";
            when "10" & x"730" => data <= x"6b";
            when "10" & x"731" => data <= x"20";
            when "10" & x"732" => data <= x"6c";
            when "10" & x"733" => data <= x"65";
            when "10" & x"734" => data <= x"6e";
            when "10" & x"735" => data <= x"20";
            when "10" & x"736" => data <= x"65";
            when "10" & x"737" => data <= x"72";
            when "10" & x"738" => data <= x"72";
            when "10" & x"739" => data <= x"6f";
            when "10" & x"73a" => data <= x"72";
            when "10" & x"73b" => data <= x"20";
            when "10" & x"73c" => data <= x"00";
            when "10" & x"73d" => data <= x"a9";
            when "10" & x"73e" => data <= x"51";
            when "10" & x"73f" => data <= x"20";
            when "10" & x"740" => data <= x"6f";
            when "10" & x"741" => data <= x"a5";
            when "10" & x"742" => data <= x"60";
            when "10" & x"743" => data <= x"20";
            when "10" & x"744" => data <= x"21";
            when "10" & x"745" => data <= x"aa";
            when "10" & x"746" => data <= x"20";
            when "10" & x"747" => data <= x"32";
            when "10" & x"748" => data <= x"a3";
            when "10" & x"749" => data <= x"d0";
            when "10" & x"74a" => data <= x"07";
            when "10" & x"74b" => data <= x"20";
            when "10" & x"74c" => data <= x"a1";
            when "10" & x"74d" => data <= x"a3";
            when "10" & x"74e" => data <= x"20";
            when "10" & x"74f" => data <= x"83";
            when "10" & x"750" => data <= x"aa";
            when "10" & x"751" => data <= x"60";
            when "10" & x"752" => data <= x"20";
            when "10" & x"753" => data <= x"1f";
            when "10" & x"754" => data <= x"a0";
            when "10" & x"755" => data <= x"c5";
            when "10" & x"756" => data <= x"4d";
            when "10" & x"757" => data <= x"4d";
            when "10" & x"758" => data <= x"43";
            when "10" & x"759" => data <= x"20";
            when "10" & x"75a" => data <= x"52";
            when "10" & x"75b" => data <= x"65";
            when "10" & x"75c" => data <= x"61";
            when "10" & x"75d" => data <= x"64";
            when "10" & x"75e" => data <= x"20";
            when "10" & x"75f" => data <= x"66";
            when "10" & x"760" => data <= x"61";
            when "10" & x"761" => data <= x"75";
            when "10" & x"762" => data <= x"6c";
            when "10" & x"763" => data <= x"74";
            when "10" & x"764" => data <= x"20";
            when "10" & x"765" => data <= x"00";
            when "10" & x"766" => data <= x"20";
            when "10" & x"767" => data <= x"21";
            when "10" & x"768" => data <= x"aa";
            when "10" & x"769" => data <= x"20";
            when "10" & x"76a" => data <= x"32";
            when "10" & x"76b" => data <= x"a3";
            when "10" & x"76c" => data <= x"d0";
            when "10" & x"76d" => data <= x"07";
            when "10" & x"76e" => data <= x"20";
            when "10" & x"76f" => data <= x"92";
            when "10" & x"770" => data <= x"a4";
            when "10" & x"771" => data <= x"20";
            when "10" & x"772" => data <= x"83";
            when "10" & x"773" => data <= x"aa";
            when "10" & x"774" => data <= x"60";
            when "10" & x"775" => data <= x"20";
            when "10" & x"776" => data <= x"1f";
            when "10" & x"777" => data <= x"a0";
            when "10" & x"778" => data <= x"c5";
            when "10" & x"779" => data <= x"4d";
            when "10" & x"77a" => data <= x"4d";
            when "10" & x"77b" => data <= x"43";
            when "10" & x"77c" => data <= x"20";
            when "10" & x"77d" => data <= x"57";
            when "10" & x"77e" => data <= x"72";
            when "10" & x"77f" => data <= x"69";
            when "10" & x"780" => data <= x"74";
            when "10" & x"781" => data <= x"65";
            when "10" & x"782" => data <= x"20";
            when "10" & x"783" => data <= x"66";
            when "10" & x"784" => data <= x"61";
            when "10" & x"785" => data <= x"75";
            when "10" & x"786" => data <= x"6c";
            when "10" & x"787" => data <= x"74";
            when "10" & x"788" => data <= x"20";
            when "10" & x"789" => data <= x"00";
            when "10" & x"78a" => data <= x"20";
            when "10" & x"78b" => data <= x"76";
            when "10" & x"78c" => data <= x"a1";
            when "10" & x"78d" => data <= x"a9";
            when "10" & x"78e" => data <= x"00";
            when "10" & x"78f" => data <= x"8d";
            when "10" & x"790" => data <= x"d6";
            when "10" & x"791" => data <= x"10";
            when "10" & x"792" => data <= x"85";
            when "10" & x"793" => data <= x"a0";
            when "10" & x"794" => data <= x"a9";
            when "10" & x"795" => data <= x"0e";
            when "10" & x"796" => data <= x"85";
            when "10" & x"797" => data <= x"a1";
            when "10" & x"798" => data <= x"60";
            when "10" & x"799" => data <= x"20";
            when "10" & x"79a" => data <= x"8a";
            when "10" & x"79b" => data <= x"a7";
            when "10" & x"79c" => data <= x"20";
            when "10" & x"79d" => data <= x"3d";
            when "10" & x"79e" => data <= x"a7";
            when "10" & x"79f" => data <= x"20";
            when "10" & x"7a0" => data <= x"43";
            when "10" & x"7a1" => data <= x"a7";
            when "10" & x"7a2" => data <= x"20";
            when "10" & x"7a3" => data <= x"be";
            when "10" & x"7a4" => data <= x"a3";
            when "10" & x"7a5" => data <= x"e6";
            when "10" & x"7a6" => data <= x"a1";
            when "10" & x"7a7" => data <= x"20";
            when "10" & x"7a8" => data <= x"be";
            when "10" & x"7a9" => data <= x"a3";
            when "10" & x"7aa" => data <= x"a0";
            when "10" & x"7ab" => data <= x"02";
            when "10" & x"7ac" => data <= x"20";
            when "10" & x"7ad" => data <= x"da";
            when "10" & x"7ae" => data <= x"a2";
            when "10" & x"7af" => data <= x"4c";
            when "10" & x"7b0" => data <= x"80";
            when "10" & x"7b1" => data <= x"a1";
            when "10" & x"7b2" => data <= x"20";
            when "10" & x"7b3" => data <= x"8a";
            when "10" & x"7b4" => data <= x"a7";
            when "10" & x"7b5" => data <= x"a9";
            when "10" & x"7b6" => data <= x"58";
            when "10" & x"7b7" => data <= x"20";
            when "10" & x"7b8" => data <= x"3f";
            when "10" & x"7b9" => data <= x"a7";
            when "10" & x"7ba" => data <= x"20";
            when "10" & x"7bb" => data <= x"66";
            when "10" & x"7bc" => data <= x"a7";
            when "10" & x"7bd" => data <= x"20";
            when "10" & x"7be" => data <= x"15";
            when "10" & x"7bf" => data <= x"a5";
            when "10" & x"7c0" => data <= x"e6";
            when "10" & x"7c1" => data <= x"a1";
            when "10" & x"7c2" => data <= x"20";
            when "10" & x"7c3" => data <= x"15";
            when "10" & x"7c4" => data <= x"a5";
            when "10" & x"7c5" => data <= x"20";
            when "10" & x"7c6" => data <= x"b4";
            when "10" & x"7c7" => data <= x"a4";
            when "10" & x"7c8" => data <= x"4c";
            when "10" & x"7c9" => data <= x"80";
            when "10" & x"7ca" => data <= x"a1";
            when "10" & x"7cb" => data <= x"60";
            when "10" & x"7cc" => data <= x"20";
            when "10" & x"7cd" => data <= x"76";
            when "10" & x"7ce" => data <= x"a1";
            when "10" & x"7cf" => data <= x"20";
            when "10" & x"7d0" => data <= x"d5";
            when "10" & x"7d1" => data <= x"a7";
            when "10" & x"7d2" => data <= x"4c";
            when "10" & x"7d3" => data <= x"80";
            when "10" & x"7d4" => data <= x"a1";
            when "10" & x"7d5" => data <= x"ae";
            when "10" & x"7d6" => data <= x"27";
            when "10" & x"7d7" => data <= x"0d";
            when "10" & x"7d8" => data <= x"f0";
            when "10" & x"7d9" => data <= x"f1";
            when "10" & x"7da" => data <= x"a9";
            when "10" & x"7db" => data <= x"01";
            when "10" & x"7dc" => data <= x"20";
            when "10" & x"7dd" => data <= x"98";
            when "10" & x"7de" => data <= x"a0";
            when "10" & x"7df" => data <= x"ae";
            when "10" & x"7e0" => data <= x"27";
            when "10" & x"7e1" => data <= x"0d";
            when "10" & x"7e2" => data <= x"2c";
            when "10" & x"7e3" => data <= x"28";
            when "10" & x"7e4" => data <= x"0d";
            when "10" & x"7e5" => data <= x"10";
            when "10" & x"7e6" => data <= x"01";
            when "10" & x"7e7" => data <= x"e8";
            when "10" & x"7e8" => data <= x"8e";
            when "10" & x"7e9" => data <= x"27";
            when "10" & x"7ea" => data <= x"0d";
            when "10" & x"7eb" => data <= x"20";
            when "10" & x"7ec" => data <= x"3d";
            when "10" & x"7ed" => data <= x"a7";
            when "10" & x"7ee" => data <= x"ae";
            when "10" & x"7ef" => data <= x"27";
            when "10" & x"7f0" => data <= x"0d";
            when "10" & x"7f1" => data <= x"e0";
            when "10" & x"7f2" => data <= x"03";
            when "10" & x"7f3" => data <= x"b0";
            when "10" & x"7f4" => data <= x"09";
            when "10" & x"7f5" => data <= x"ad";
            when "10" & x"7f6" => data <= x"29";
            when "10" & x"7f7" => data <= x"0d";
            when "10" & x"7f8" => data <= x"d0";
            when "10" & x"7f9" => data <= x"46";
            when "10" & x"7fa" => data <= x"e0";
            when "10" & x"7fb" => data <= x"01";
            when "10" & x"7fc" => data <= x"f0";
            when "10" & x"7fd" => data <= x"39";
            when "10" & x"7fe" => data <= x"2c";
            when "10" & x"7ff" => data <= x"28";
            when "10" & x"800" => data <= x"0d";
            when "10" & x"801" => data <= x"10";
            when "10" & x"802" => data <= x"0e";
            when "10" & x"803" => data <= x"20";
            when "10" & x"804" => data <= x"43";
            when "10" & x"805" => data <= x"a7";
            when "10" & x"806" => data <= x"a0";
            when "10" & x"807" => data <= x"00";
            when "10" & x"808" => data <= x"8c";
            when "10" & x"809" => data <= x"28";
            when "10" & x"80a" => data <= x"0d";
            when "10" & x"80b" => data <= x"20";
            when "10" & x"80c" => data <= x"da";
            when "10" & x"80d" => data <= x"a2";
            when "10" & x"80e" => data <= x"4c";
            when "10" & x"80f" => data <= x"19";
            when "10" & x"810" => data <= x"a8";
            when "10" & x"811" => data <= x"20";
            when "10" & x"812" => data <= x"43";
            when "10" & x"813" => data <= x"a7";
            when "10" & x"814" => data <= x"20";
            when "10" & x"815" => data <= x"be";
            when "10" & x"816" => data <= x"a3";
            when "10" & x"817" => data <= x"e6";
            when "10" & x"818" => data <= x"a1";
            when "10" & x"819" => data <= x"20";
            when "10" & x"81a" => data <= x"be";
            when "10" & x"81b" => data <= x"a3";
            when "10" & x"81c" => data <= x"e6";
            when "10" & x"81d" => data <= x"a1";
            when "10" & x"81e" => data <= x"a0";
            when "10" & x"81f" => data <= x"02";
            when "10" & x"820" => data <= x"20";
            when "10" & x"821" => data <= x"da";
            when "10" & x"822" => data <= x"a2";
            when "10" & x"823" => data <= x"20";
            when "10" & x"824" => data <= x"61";
            when "10" & x"825" => data <= x"aa";
            when "10" & x"826" => data <= x"ae";
            when "10" & x"827" => data <= x"27";
            when "10" & x"828" => data <= x"0d";
            when "10" & x"829" => data <= x"ca";
            when "10" & x"82a" => data <= x"ca";
            when "10" & x"82b" => data <= x"f0";
            when "10" & x"82c" => data <= x"9e";
            when "10" & x"82d" => data <= x"8e";
            when "10" & x"82e" => data <= x"27";
            when "10" & x"82f" => data <= x"0d";
            when "10" & x"830" => data <= x"e0";
            when "10" & x"831" => data <= x"03";
            when "10" & x"832" => data <= x"b0";
            when "10" & x"833" => data <= x"dd";
            when "10" & x"834" => data <= x"4c";
            when "10" & x"835" => data <= x"f5";
            when "10" & x"836" => data <= x"a7";
            when "10" & x"837" => data <= x"20";
            when "10" & x"838" => data <= x"43";
            when "10" & x"839" => data <= x"a7";
            when "10" & x"83a" => data <= x"20";
            when "10" & x"83b" => data <= x"be";
            when "10" & x"83c" => data <= x"a3";
            when "10" & x"83d" => data <= x"4c";
            when "10" & x"83e" => data <= x"6d";
            when "10" & x"83f" => data <= x"a8";
            when "10" & x"840" => data <= x"20";
            when "10" & x"841" => data <= x"43";
            when "10" & x"842" => data <= x"a7";
            when "10" & x"843" => data <= x"2c";
            when "10" & x"844" => data <= x"28";
            when "10" & x"845" => data <= x"0d";
            when "10" & x"846" => data <= x"10";
            when "10" & x"847" => data <= x"0b";
            when "10" & x"848" => data <= x"a0";
            when "10" & x"849" => data <= x"00";
            when "10" & x"84a" => data <= x"8c";
            when "10" & x"84b" => data <= x"28";
            when "10" & x"84c" => data <= x"0d";
            when "10" & x"84d" => data <= x"20";
            when "10" & x"84e" => data <= x"da";
            when "10" & x"84f" => data <= x"a2";
            when "10" & x"850" => data <= x"4c";
            when "10" & x"851" => data <= x"5d";
            when "10" & x"852" => data <= x"a8";
            when "10" & x"853" => data <= x"ce";
            when "10" & x"854" => data <= x"27";
            when "10" & x"855" => data <= x"0d";
            when "10" & x"856" => data <= x"f0";
            when "10" & x"857" => data <= x"05";
            when "10" & x"858" => data <= x"20";
            when "10" & x"859" => data <= x"be";
            when "10" & x"85a" => data <= x"a3";
            when "10" & x"85b" => data <= x"e6";
            when "10" & x"85c" => data <= x"a1";
            when "10" & x"85d" => data <= x"20";
            when "10" & x"85e" => data <= x"f5";
            when "10" & x"85f" => data <= x"a3";
            when "10" & x"860" => data <= x"98";
            when "10" & x"861" => data <= x"49";
            when "10" & x"862" => data <= x"ff";
            when "10" & x"863" => data <= x"a8";
            when "10" & x"864" => data <= x"c8";
            when "10" & x"865" => data <= x"20";
            when "10" & x"866" => data <= x"da";
            when "10" & x"867" => data <= x"a2";
            when "10" & x"868" => data <= x"ad";
            when "10" & x"869" => data <= x"27";
            when "10" & x"86a" => data <= x"0d";
            when "10" & x"86b" => data <= x"d0";
            when "10" & x"86c" => data <= x"05";
            when "10" & x"86d" => data <= x"a0";
            when "10" & x"86e" => data <= x"00";
            when "10" & x"86f" => data <= x"20";
            when "10" & x"870" => data <= x"da";
            when "10" & x"871" => data <= x"a2";
            when "10" & x"872" => data <= x"a0";
            when "10" & x"873" => data <= x"02";
            when "10" & x"874" => data <= x"4c";
            when "10" & x"875" => data <= x"da";
            when "10" & x"876" => data <= x"a2";
            when "10" & x"877" => data <= x"60";
            when "10" & x"878" => data <= x"20";
            when "10" & x"879" => data <= x"76";
            when "10" & x"87a" => data <= x"a1";
            when "10" & x"87b" => data <= x"20";
            when "10" & x"87c" => data <= x"81";
            when "10" & x"87d" => data <= x"a8";
            when "10" & x"87e" => data <= x"4c";
            when "10" & x"87f" => data <= x"80";
            when "10" & x"880" => data <= x"a1";
            when "10" & x"881" => data <= x"ae";
            when "10" & x"882" => data <= x"27";
            when "10" & x"883" => data <= x"0d";
            when "10" & x"884" => data <= x"f0";
            when "10" & x"885" => data <= x"f1";
            when "10" & x"886" => data <= x"a9";
            when "10" & x"887" => data <= x"00";
            when "10" & x"888" => data <= x"20";
            when "10" & x"889" => data <= x"98";
            when "10" & x"88a" => data <= x"a0";
            when "10" & x"88b" => data <= x"a9";
            when "10" & x"88c" => data <= x"58";
            when "10" & x"88d" => data <= x"20";
            when "10" & x"88e" => data <= x"3f";
            when "10" & x"88f" => data <= x"a7";
            when "10" & x"890" => data <= x"ae";
            when "10" & x"891" => data <= x"27";
            when "10" & x"892" => data <= x"0d";
            when "10" & x"893" => data <= x"2c";
            when "10" & x"894" => data <= x"28";
            when "10" & x"895" => data <= x"0d";
            when "10" & x"896" => data <= x"10";
            when "10" & x"897" => data <= x"3a";
            when "10" & x"898" => data <= x"a9";
            when "10" & x"899" => data <= x"00";
            when "10" & x"89a" => data <= x"8d";
            when "10" & x"89b" => data <= x"28";
            when "10" & x"89c" => data <= x"0d";
            when "10" & x"89d" => data <= x"a9";
            when "10" & x"89e" => data <= x"ff";
            when "10" & x"89f" => data <= x"8d";
            when "10" & x"8a0" => data <= x"82";
            when "10" & x"8a1" => data <= x"10";
            when "10" & x"8a2" => data <= x"a9";
            when "10" & x"8a3" => data <= x"51";
            when "10" & x"8a4" => data <= x"8d";
            when "10" & x"8a5" => data <= x"43";
            when "10" & x"8a6" => data <= x"0d";
            when "10" & x"8a7" => data <= x"20";
            when "10" & x"8a8" => data <= x"43";
            when "10" & x"8a9" => data <= x"a7";
            when "10" & x"8aa" => data <= x"20";
            when "10" & x"8ab" => data <= x"62";
            when "10" & x"8ac" => data <= x"a4";
            when "10" & x"8ad" => data <= x"a0";
            when "10" & x"8ae" => data <= x"00";
            when "10" & x"8af" => data <= x"20";
            when "10" & x"8b0" => data <= x"da";
            when "10" & x"8b1" => data <= x"a2";
            when "10" & x"8b2" => data <= x"a0";
            when "10" & x"8b3" => data <= x"02";
            when "10" & x"8b4" => data <= x"20";
            when "10" & x"8b5" => data <= x"da";
            when "10" & x"8b6" => data <= x"a2";
            when "10" & x"8b7" => data <= x"a9";
            when "10" & x"8b8" => data <= x"58";
            when "10" & x"8b9" => data <= x"8d";
            when "10" & x"8ba" => data <= x"43";
            when "10" & x"8bb" => data <= x"0d";
            when "10" & x"8bc" => data <= x"20";
            when "10" & x"8bd" => data <= x"66";
            when "10" & x"8be" => data <= x"a7";
            when "10" & x"8bf" => data <= x"20";
            when "10" & x"8c0" => data <= x"51";
            when "10" & x"8c1" => data <= x"a5";
            when "10" & x"8c2" => data <= x"20";
            when "10" & x"8c3" => data <= x"15";
            when "10" & x"8c4" => data <= x"a5";
            when "10" & x"8c5" => data <= x"20";
            when "10" & x"8c6" => data <= x"b4";
            when "10" & x"8c7" => data <= x"a4";
            when "10" & x"8c8" => data <= x"ce";
            when "10" & x"8c9" => data <= x"27";
            when "10" & x"8ca" => data <= x"0d";
            when "10" & x"8cb" => data <= x"f0";
            when "10" & x"8cc" => data <= x"aa";
            when "10" & x"8cd" => data <= x"e6";
            when "10" & x"8ce" => data <= x"a1";
            when "10" & x"8cf" => data <= x"20";
            when "10" & x"8d0" => data <= x"61";
            when "10" & x"8d1" => data <= x"aa";
            when "10" & x"8d2" => data <= x"ae";
            when "10" & x"8d3" => data <= x"27";
            when "10" & x"8d4" => data <= x"0d";
            when "10" & x"8d5" => data <= x"f0";
            when "10" & x"8d6" => data <= x"46";
            when "10" & x"8d7" => data <= x"ca";
            when "10" & x"8d8" => data <= x"d0";
            when "10" & x"8d9" => data <= x"2b";
            when "10" & x"8da" => data <= x"a9";
            when "10" & x"8db" => data <= x"ff";
            when "10" & x"8dc" => data <= x"8d";
            when "10" & x"8dd" => data <= x"82";
            when "10" & x"8de" => data <= x"10";
            when "10" & x"8df" => data <= x"a9";
            when "10" & x"8e0" => data <= x"51";
            when "10" & x"8e1" => data <= x"8d";
            when "10" & x"8e2" => data <= x"43";
            when "10" & x"8e3" => data <= x"0d";
            when "10" & x"8e4" => data <= x"20";
            when "10" & x"8e5" => data <= x"43";
            when "10" & x"8e6" => data <= x"a7";
            when "10" & x"8e7" => data <= x"a0";
            when "10" & x"8e8" => data <= x"00";
            when "10" & x"8e9" => data <= x"20";
            when "10" & x"8ea" => data <= x"da";
            when "10" & x"8eb" => data <= x"a2";
            when "10" & x"8ec" => data <= x"20";
            when "10" & x"8ed" => data <= x"62";
            when "10" & x"8ee" => data <= x"a4";
            when "10" & x"8ef" => data <= x"a0";
            when "10" & x"8f0" => data <= x"02";
            when "10" & x"8f1" => data <= x"20";
            when "10" & x"8f2" => data <= x"da";
            when "10" & x"8f3" => data <= x"a2";
            when "10" & x"8f4" => data <= x"a9";
            when "10" & x"8f5" => data <= x"58";
            when "10" & x"8f6" => data <= x"8d";
            when "10" & x"8f7" => data <= x"43";
            when "10" & x"8f8" => data <= x"0d";
            when "10" & x"8f9" => data <= x"20";
            when "10" & x"8fa" => data <= x"66";
            when "10" & x"8fb" => data <= x"a7";
            when "10" & x"8fc" => data <= x"20";
            when "10" & x"8fd" => data <= x"15";
            when "10" & x"8fe" => data <= x"a5";
            when "10" & x"8ff" => data <= x"20";
            when "10" & x"900" => data <= x"51";
            when "10" & x"901" => data <= x"a5";
            when "10" & x"902" => data <= x"4c";
            when "10" & x"903" => data <= x"b4";
            when "10" & x"904" => data <= x"a4";
            when "10" & x"905" => data <= x"20";
            when "10" & x"906" => data <= x"66";
            when "10" & x"907" => data <= x"a7";
            when "10" & x"908" => data <= x"20";
            when "10" & x"909" => data <= x"15";
            when "10" & x"90a" => data <= x"a5";
            when "10" & x"90b" => data <= x"e6";
            when "10" & x"90c" => data <= x"a1";
            when "10" & x"90d" => data <= x"20";
            when "10" & x"90e" => data <= x"15";
            when "10" & x"90f" => data <= x"a5";
            when "10" & x"910" => data <= x"e6";
            when "10" & x"911" => data <= x"a1";
            when "10" & x"912" => data <= x"20";
            when "10" & x"913" => data <= x"b4";
            when "10" & x"914" => data <= x"a4";
            when "10" & x"915" => data <= x"ce";
            when "10" & x"916" => data <= x"27";
            when "10" & x"917" => data <= x"0d";
            when "10" & x"918" => data <= x"ce";
            when "10" & x"919" => data <= x"27";
            when "10" & x"91a" => data <= x"0d";
            when "10" & x"91b" => data <= x"d0";
            when "10" & x"91c" => data <= x"b2";
            when "10" & x"91d" => data <= x"60";
            when "10" & x"91e" => data <= x"a9";
            when "10" & x"91f" => data <= x"51";
            when "10" & x"920" => data <= x"20";
            when "10" & x"921" => data <= x"6f";
            when "10" & x"922" => data <= x"a5";
            when "10" & x"923" => data <= x"60";
            when "10" & x"924" => data <= x"20";
            when "10" & x"925" => data <= x"76";
            when "10" & x"926" => data <= x"a1";
            when "10" & x"927" => data <= x"20";
            when "10" & x"928" => data <= x"43";
            when "10" & x"929" => data <= x"a7";
            when "10" & x"92a" => data <= x"a9";
            when "10" & x"92b" => data <= x"5f";
            when "10" & x"92c" => data <= x"85";
            when "10" & x"92d" => data <= x"a0";
            when "10" & x"92e" => data <= x"a9";
            when "10" & x"92f" => data <= x"0d";
            when "10" & x"930" => data <= x"85";
            when "10" & x"931" => data <= x"a1";
            when "10" & x"932" => data <= x"a9";
            when "10" & x"933" => data <= x"08";
            when "10" & x"934" => data <= x"8d";
            when "10" & x"935" => data <= x"29";
            when "10" & x"936" => data <= x"0d";
            when "10" & x"937" => data <= x"20";
            when "10" & x"938" => data <= x"f5";
            when "10" & x"939" => data <= x"a3";
            when "10" & x"93a" => data <= x"a0";
            when "10" & x"93b" => data <= x"f8";
            when "10" & x"93c" => data <= x"20";
            when "10" & x"93d" => data <= x"da";
            when "10" & x"93e" => data <= x"a2";
            when "10" & x"93f" => data <= x"a9";
            when "10" & x"940" => data <= x"67";
            when "10" & x"941" => data <= x"85";
            when "10" & x"942" => data <= x"a0";
            when "10" & x"943" => data <= x"a9";
            when "10" & x"944" => data <= x"08";
            when "10" & x"945" => data <= x"8d";
            when "10" & x"946" => data <= x"29";
            when "10" & x"947" => data <= x"0d";
            when "10" & x"948" => data <= x"20";
            when "10" & x"949" => data <= x"f5";
            when "10" & x"94a" => data <= x"a3";
            when "10" & x"94b" => data <= x"a0";
            when "10" & x"94c" => data <= x"fa";
            when "10" & x"94d" => data <= x"20";
            when "10" & x"94e" => data <= x"da";
            when "10" & x"94f" => data <= x"a2";
            when "10" & x"950" => data <= x"ad";
            when "10" & x"951" => data <= x"4f";
            when "10" & x"952" => data <= x"0d";
            when "10" & x"953" => data <= x"c9";
            when "10" & x"954" => data <= x"02";
            when "10" & x"955" => data <= x"f0";
            when "10" & x"956" => data <= x"1e";
            when "10" & x"957" => data <= x"18";
            when "10" & x"958" => data <= x"ad";
            when "10" & x"959" => data <= x"47";
            when "10" & x"95a" => data <= x"0d";
            when "10" & x"95b" => data <= x"69";
            when "10" & x"95c" => data <= x"90";
            when "10" & x"95d" => data <= x"8d";
            when "10" & x"95e" => data <= x"47";
            when "10" & x"95f" => data <= x"0d";
            when "10" & x"960" => data <= x"ad";
            when "10" & x"961" => data <= x"46";
            when "10" & x"962" => data <= x"0d";
            when "10" & x"963" => data <= x"69";
            when "10" & x"964" => data <= x"01";
            when "10" & x"965" => data <= x"8d";
            when "10" & x"966" => data <= x"46";
            when "10" & x"967" => data <= x"0d";
            when "10" & x"968" => data <= x"90";
            when "10" & x"969" => data <= x"08";
            when "10" & x"96a" => data <= x"ee";
            when "10" & x"96b" => data <= x"45";
            when "10" & x"96c" => data <= x"0d";
            when "10" & x"96d" => data <= x"f0";
            when "10" & x"96e" => data <= x"03";
            when "10" & x"96f" => data <= x"ee";
            when "10" & x"970" => data <= x"44";
            when "10" & x"971" => data <= x"0d";
            when "10" & x"972" => data <= x"4c";
            when "10" & x"973" => data <= x"8b";
            when "10" & x"974" => data <= x"a9";
            when "10" & x"975" => data <= x"18";
            when "10" & x"976" => data <= x"ad";
            when "10" & x"977" => data <= x"46";
            when "10" & x"978" => data <= x"0d";
            when "10" & x"979" => data <= x"69";
            when "10" & x"97a" => data <= x"20";
            when "10" & x"97b" => data <= x"8d";
            when "10" & x"97c" => data <= x"46";
            when "10" & x"97d" => data <= x"0d";
            when "10" & x"97e" => data <= x"ad";
            when "10" & x"97f" => data <= x"45";
            when "10" & x"980" => data <= x"0d";
            when "10" & x"981" => data <= x"69";
            when "10" & x"982" => data <= x"03";
            when "10" & x"983" => data <= x"8d";
            when "10" & x"984" => data <= x"45";
            when "10" & x"985" => data <= x"0d";
            when "10" & x"986" => data <= x"90";
            when "10" & x"987" => data <= x"03";
            when "10" & x"988" => data <= x"ee";
            when "10" & x"989" => data <= x"44";
            when "10" & x"98a" => data <= x"0d";
            when "10" & x"98b" => data <= x"4c";
            when "10" & x"98c" => data <= x"80";
            when "10" & x"98d" => data <= x"a1";
            when "10" & x"98e" => data <= x"60";
            when "10" & x"98f" => data <= x"a9";
            when "10" & x"990" => data <= x"00";
            when "10" & x"991" => data <= x"8d";
            when "10" & x"992" => data <= x"50";
            when "10" & x"993" => data <= x"0d";
            when "10" & x"994" => data <= x"8d";
            when "10" & x"995" => data <= x"51";
            when "10" & x"996" => data <= x"0d";
            when "10" & x"997" => data <= x"20";
            when "10" & x"998" => data <= x"eb";
            when "10" & x"999" => data <= x"a9";
            when "10" & x"99a" => data <= x"a9";
            when "10" & x"99b" => data <= x"7a";
            when "10" & x"99c" => data <= x"20";
            when "10" & x"99d" => data <= x"f4";
            when "10" & x"99e" => data <= x"ff";
            when "10" & x"99f" => data <= x"8a";
            when "10" & x"9a0" => data <= x"30";
            when "10" & x"9a1" => data <= x"0d";
            when "10" & x"9a2" => data <= x"c9";
            when "10" & x"9a3" => data <= x"51";
            when "10" & x"9a4" => data <= x"f0";
            when "10" & x"9a5" => data <= x"04";
            when "10" & x"9a6" => data <= x"c9";
            when "10" & x"9a7" => data <= x"42";
            when "10" & x"9a8" => data <= x"d0";
            when "10" & x"9a9" => data <= x"e4";
            when "10" & x"9aa" => data <= x"a9";
            when "10" & x"9ab" => data <= x"78";
            when "10" & x"9ac" => data <= x"20";
            when "10" & x"9ad" => data <= x"f4";
            when "10" & x"9ae" => data <= x"ff";
            when "10" & x"9af" => data <= x"8e";
            when "10" & x"9b0" => data <= x"52";
            when "10" & x"9b1" => data <= x"0d";
            when "10" & x"9b2" => data <= x"4c";
            when "10" & x"9b3" => data <= x"20";
            when "10" & x"9b4" => data <= x"93";
            when "10" & x"9b5" => data <= x"ae";
            when "10" & x"9b6" => data <= x"4a";
            when "10" & x"9b7" => data <= x"0d";
            when "10" & x"9b8" => data <= x"18";
            when "10" & x"9b9" => data <= x"a9";
            when "10" & x"9ba" => data <= x"80";
            when "10" & x"9bb" => data <= x"2a";
            when "10" & x"9bc" => data <= x"2a";
            when "10" & x"9bd" => data <= x"ca";
            when "10" & x"9be" => data <= x"d0";
            when "10" & x"9bf" => data <= x"fb";
            when "10" & x"9c0" => data <= x"8d";
            when "10" & x"9c1" => data <= x"4b";
            when "10" & x"9c2" => data <= x"0d";
            when "10" & x"9c3" => data <= x"0a";
            when "10" & x"9c4" => data <= x"8d";
            when "10" & x"9c5" => data <= x"4e";
            when "10" & x"9c6" => data <= x"0d";
            when "10" & x"9c7" => data <= x"aa";
            when "10" & x"9c8" => data <= x"18";
            when "10" & x"9c9" => data <= x"6d";
            when "10" & x"9ca" => data <= x"4b";
            when "10" & x"9cb" => data <= x"0d";
            when "10" & x"9cc" => data <= x"8d";
            when "10" & x"9cd" => data <= x"4c";
            when "10" & x"9ce" => data <= x"0d";
            when "10" & x"9cf" => data <= x"8a";
            when "10" & x"9d0" => data <= x"49";
            when "10" & x"9d1" => data <= x"ff";
            when "10" & x"9d2" => data <= x"8d";
            when "10" & x"9d3" => data <= x"4d";
            when "10" & x"9d4" => data <= x"0d";
            when "10" & x"9d5" => data <= x"60";
            when "10" & x"9d6" => data <= x"ad";
            when "10" & x"9d7" => data <= x"b2";
            when "10" & x"9d8" => data <= x"fc";
            when "10" & x"9d9" => data <= x"8d";
            when "10" & x"9da" => data <= x"50";
            when "10" & x"9db" => data <= x"0d";
            when "10" & x"9dc" => data <= x"49";
            when "10" & x"9dd" => data <= x"ff";
            when "10" & x"9de" => data <= x"8d";
            when "10" & x"9df" => data <= x"51";
            when "10" & x"9e0" => data <= x"0d";
            when "10" & x"9e1" => data <= x"ad";
            when "10" & x"9e2" => data <= x"b0";
            when "10" & x"9e3" => data <= x"fc";
            when "10" & x"9e4" => data <= x"4d";
            when "10" & x"9e5" => data <= x"51";
            when "10" & x"9e6" => data <= x"0d";
            when "10" & x"9e7" => data <= x"8d";
            when "10" & x"9e8" => data <= x"51";
            when "10" & x"9e9" => data <= x"0d";
            when "10" & x"9ea" => data <= x"60";
            when "10" & x"9eb" => data <= x"a9";
            when "10" & x"9ec" => data <= x"00";
            when "10" & x"9ed" => data <= x"8d";
            when "10" & x"9ee" => data <= x"3f";
            when "10" & x"9ef" => data <= x"0d";
            when "10" & x"9f0" => data <= x"8d";
            when "10" & x"9f1" => data <= x"4f";
            when "10" & x"9f2" => data <= x"0d";
            when "10" & x"9f3" => data <= x"a2";
            when "10" & x"9f4" => data <= x"04";
            when "10" & x"9f5" => data <= x"8e";
            when "10" & x"9f6" => data <= x"4a";
            when "10" & x"9f7" => data <= x"0d";
            when "10" & x"9f8" => data <= x"20";
            when "10" & x"9f9" => data <= x"b5";
            when "10" & x"9fa" => data <= x"a9";
            when "10" & x"9fb" => data <= x"20";
            when "10" & x"9fc" => data <= x"43";
            when "10" & x"9fd" => data <= x"a6";
            when "10" & x"9fe" => data <= x"c9";
            when "10" & x"9ff" => data <= x"ff";
            when "10" & x"a00" => data <= x"f0";
            when "10" & x"a01" => data <= x"1e";
            when "10" & x"a02" => data <= x"ae";
            when "10" & x"a03" => data <= x"4a";
            when "10" & x"a04" => data <= x"0d";
            when "10" & x"a05" => data <= x"ca";
            when "10" & x"a06" => data <= x"d0";
            when "10" & x"a07" => data <= x"ed";
            when "10" & x"a08" => data <= x"8e";
            when "10" & x"a09" => data <= x"4a";
            when "10" & x"a0a" => data <= x"0d";
            when "10" & x"a0b" => data <= x"8e";
            when "10" & x"a0c" => data <= x"4f";
            when "10" & x"a0d" => data <= x"0d";
            when "10" & x"a0e" => data <= x"ad";
            when "10" & x"a0f" => data <= x"3f";
            when "10" & x"a10" => data <= x"0d";
            when "10" & x"a11" => data <= x"d0";
            when "10" & x"a12" => data <= x"0a";
            when "10" & x"a13" => data <= x"a2";
            when "10" & x"a14" => data <= x"08";
            when "10" & x"a15" => data <= x"8e";
            when "10" & x"a16" => data <= x"3f";
            when "10" & x"a17" => data <= x"0d";
            when "10" & x"a18" => data <= x"a2";
            when "10" & x"a19" => data <= x"01";
            when "10" & x"a1a" => data <= x"4c";
            when "10" & x"a1b" => data <= x"f5";
            when "10" & x"a1c" => data <= x"a9";
            when "10" & x"a1d" => data <= x"20";
            when "10" & x"a1e" => data <= x"07";
            when "10" & x"a1f" => data <= x"a7";
            when "10" & x"a20" => data <= x"60";
            when "10" & x"a21" => data <= x"ad";
            when "10" & x"a22" => data <= x"4f";
            when "10" & x"a23" => data <= x"0d";
            when "10" & x"a24" => data <= x"c9";
            when "10" & x"a25" => data <= x"02";
            when "10" & x"a26" => data <= x"d0";
            when "10" & x"a27" => data <= x"20";
            when "10" & x"a28" => data <= x"ad";
            when "10" & x"a29" => data <= x"26";
            when "10" & x"a2a" => data <= x"0d";
            when "10" & x"a2b" => data <= x"18";
            when "10" & x"a2c" => data <= x"ac";
            when "10" & x"a2d" => data <= x"25";
            when "10" & x"a2e" => data <= x"0d";
            when "10" & x"a2f" => data <= x"ae";
            when "10" & x"a30" => data <= x"24";
            when "10" & x"a31" => data <= x"0d";
            when "10" & x"a32" => data <= x"ad";
            when "10" & x"a33" => data <= x"23";
            when "10" & x"a34" => data <= x"0d";
            when "10" & x"a35" => data <= x"0a";
            when "10" & x"a36" => data <= x"8d";
            when "10" & x"a37" => data <= x"24";
            when "10" & x"a38" => data <= x"0d";
            when "10" & x"a39" => data <= x"8a";
            when "10" & x"a3a" => data <= x"2a";
            when "10" & x"a3b" => data <= x"8d";
            when "10" & x"a3c" => data <= x"25";
            when "10" & x"a3d" => data <= x"0d";
            when "10" & x"a3e" => data <= x"98";
            when "10" & x"a3f" => data <= x"2a";
            when "10" & x"a40" => data <= x"8d";
            when "10" & x"a41" => data <= x"26";
            when "10" & x"a42" => data <= x"0d";
            when "10" & x"a43" => data <= x"a9";
            when "10" & x"a44" => data <= x"00";
            when "10" & x"a45" => data <= x"8d";
            when "10" & x"a46" => data <= x"23";
            when "10" & x"a47" => data <= x"0d";
            when "10" & x"a48" => data <= x"ad";
            when "10" & x"a49" => data <= x"23";
            when "10" & x"a4a" => data <= x"0d";
            when "10" & x"a4b" => data <= x"8d";
            when "10" & x"a4c" => data <= x"47";
            when "10" & x"a4d" => data <= x"0d";
            when "10" & x"a4e" => data <= x"ad";
            when "10" & x"a4f" => data <= x"24";
            when "10" & x"a50" => data <= x"0d";
            when "10" & x"a51" => data <= x"8d";
            when "10" & x"a52" => data <= x"46";
            when "10" & x"a53" => data <= x"0d";
            when "10" & x"a54" => data <= x"ad";
            when "10" & x"a55" => data <= x"25";
            when "10" & x"a56" => data <= x"0d";
            when "10" & x"a57" => data <= x"8d";
            when "10" & x"a58" => data <= x"45";
            when "10" & x"a59" => data <= x"0d";
            when "10" & x"a5a" => data <= x"ad";
            when "10" & x"a5b" => data <= x"26";
            when "10" & x"a5c" => data <= x"0d";
            when "10" & x"a5d" => data <= x"8d";
            when "10" & x"a5e" => data <= x"44";
            when "10" & x"a5f" => data <= x"0d";
            when "10" & x"a60" => data <= x"60";
            when "10" & x"a61" => data <= x"18";
            when "10" & x"a62" => data <= x"a9";
            when "10" & x"a63" => data <= x"01";
            when "10" & x"a64" => data <= x"6d";
            when "10" & x"a65" => data <= x"23";
            when "10" & x"a66" => data <= x"0d";
            when "10" & x"a67" => data <= x"8d";
            when "10" & x"a68" => data <= x"23";
            when "10" & x"a69" => data <= x"0d";
            when "10" & x"a6a" => data <= x"ad";
            when "10" & x"a6b" => data <= x"24";
            when "10" & x"a6c" => data <= x"0d";
            when "10" & x"a6d" => data <= x"69";
            when "10" & x"a6e" => data <= x"00";
            when "10" & x"a6f" => data <= x"8d";
            when "10" & x"a70" => data <= x"24";
            when "10" & x"a71" => data <= x"0d";
            when "10" & x"a72" => data <= x"ad";
            when "10" & x"a73" => data <= x"25";
            when "10" & x"a74" => data <= x"0d";
            when "10" & x"a75" => data <= x"69";
            when "10" & x"a76" => data <= x"00";
            when "10" & x"a77" => data <= x"8d";
            when "10" & x"a78" => data <= x"25";
            when "10" & x"a79" => data <= x"0d";
            when "10" & x"a7a" => data <= x"ad";
            when "10" & x"a7b" => data <= x"26";
            when "10" & x"a7c" => data <= x"0d";
            when "10" & x"a7d" => data <= x"69";
            when "10" & x"a7e" => data <= x"00";
            when "10" & x"a7f" => data <= x"8d";
            when "10" & x"a80" => data <= x"26";
            when "10" & x"a81" => data <= x"0d";
            when "10" & x"a82" => data <= x"60";
            when "10" & x"a83" => data <= x"ad";
            when "10" & x"a84" => data <= x"4f";
            when "10" & x"a85" => data <= x"0d";
            when "10" & x"a86" => data <= x"c9";
            when "10" & x"a87" => data <= x"02";
            when "10" & x"a88" => data <= x"d0";
            when "10" & x"a89" => data <= x"1c";
            when "10" & x"a8a" => data <= x"ac";
            when "10" & x"a8b" => data <= x"24";
            when "10" & x"a8c" => data <= x"0d";
            when "10" & x"a8d" => data <= x"ae";
            when "10" & x"a8e" => data <= x"25";
            when "10" & x"a8f" => data <= x"0d";
            when "10" & x"a90" => data <= x"ad";
            when "10" & x"a91" => data <= x"26";
            when "10" & x"a92" => data <= x"0d";
            when "10" & x"a93" => data <= x"4a";
            when "10" & x"a94" => data <= x"8d";
            when "10" & x"a95" => data <= x"25";
            when "10" & x"a96" => data <= x"0d";
            when "10" & x"a97" => data <= x"8a";
            when "10" & x"a98" => data <= x"6a";
            when "10" & x"a99" => data <= x"8d";
            when "10" & x"a9a" => data <= x"24";
            when "10" & x"a9b" => data <= x"0d";
            when "10" & x"a9c" => data <= x"98";
            when "10" & x"a9d" => data <= x"6a";
            when "10" & x"a9e" => data <= x"8d";
            when "10" & x"a9f" => data <= x"23";
            when "10" & x"aa0" => data <= x"0d";
            when "10" & x"aa1" => data <= x"a9";
            when "10" & x"aa2" => data <= x"00";
            when "10" & x"aa3" => data <= x"8d";
            when "10" & x"aa4" => data <= x"26";
            when "10" & x"aa5" => data <= x"0d";
            when "10" & x"aa6" => data <= x"60";
            when "10" & x"aa7" => data <= x"ad";
            when "10" & x"aa8" => data <= x"05";
            when "10" & x"aa9" => data <= x"0d";
            when "10" & x"aaa" => data <= x"c9";
            when "10" & x"aab" => data <= x"54";
            when "10" & x"aac" => data <= x"d0";
            when "10" & x"aad" => data <= x"15";
            when "10" & x"aae" => data <= x"ad";
            when "10" & x"aaf" => data <= x"06";
            when "10" & x"ab0" => data <= x"0d";
            when "10" & x"ab1" => data <= x"4d";
            when "10" & x"ab2" => data <= x"0a";
            when "10" & x"ab3" => data <= x"0d";
            when "10" & x"ab4" => data <= x"c9";
            when "10" & x"ab5" => data <= x"ff";
            when "10" & x"ab6" => data <= x"d0";
            when "10" & x"ab7" => data <= x"0b";
            when "10" & x"ab8" => data <= x"ad";
            when "10" & x"ab9" => data <= x"07";
            when "10" & x"aba" => data <= x"0d";
            when "10" & x"abb" => data <= x"4d";
            when "10" & x"abc" => data <= x"0b";
            when "10" & x"abd" => data <= x"0d";
            when "10" & x"abe" => data <= x"c9";
            when "10" & x"abf" => data <= x"ff";
            when "10" & x"ac0" => data <= x"d0";
            when "10" & x"ac1" => data <= x"01";
            when "10" & x"ac2" => data <= x"60";
            when "10" & x"ac3" => data <= x"a2";
            when "10" & x"ac4" => data <= x"0b";
            when "10" & x"ac5" => data <= x"bd";
            when "10" & x"ac6" => data <= x"22";
            when "10" & x"ac7" => data <= x"0d";
            when "10" & x"ac8" => data <= x"48";
            when "10" & x"ac9" => data <= x"ca";
            when "10" & x"aca" => data <= x"d0";
            when "10" & x"acb" => data <= x"f9";
            when "10" & x"acc" => data <= x"a9";
            when "10" & x"acd" => data <= x"00";
            when "10" & x"ace" => data <= x"8d";
            when "10" & x"acf" => data <= x"23";
            when "10" & x"ad0" => data <= x"0d";
            when "10" & x"ad1" => data <= x"8d";
            when "10" & x"ad2" => data <= x"24";
            when "10" & x"ad3" => data <= x"0d";
            when "10" & x"ad4" => data <= x"8d";
            when "10" & x"ad5" => data <= x"25";
            when "10" & x"ad6" => data <= x"0d";
            when "10" & x"ad7" => data <= x"8d";
            when "10" & x"ad8" => data <= x"26";
            when "10" & x"ad9" => data <= x"0d";
            when "10" & x"ada" => data <= x"20";
            when "10" & x"adb" => data <= x"99";
            when "10" & x"adc" => data <= x"a7";
            when "10" & x"add" => data <= x"a9";
            when "10" & x"ade" => data <= x"dd";
            when "10" & x"adf" => data <= x"8d";
            when "10" & x"ae0" => data <= x"82";
            when "10" & x"ae1" => data <= x"10";
            when "10" & x"ae2" => data <= x"20";
            when "10" & x"ae3" => data <= x"00";
            when "10" & x"ae4" => data <= x"ab";
            when "10" & x"ae5" => data <= x"f0";
            when "10" & x"ae6" => data <= x"29";
            when "10" & x"ae7" => data <= x"a9";
            when "10" & x"ae8" => data <= x"00";
            when "10" & x"ae9" => data <= x"8d";
            when "10" & x"aea" => data <= x"06";
            when "10" & x"aeb" => data <= x"0d";
            when "10" & x"aec" => data <= x"8d";
            when "10" & x"aed" => data <= x"07";
            when "10" & x"aee" => data <= x"0d";
            when "10" & x"aef" => data <= x"8d";
            when "10" & x"af0" => data <= x"08";
            when "10" & x"af1" => data <= x"0d";
            when "10" & x"af2" => data <= x"8d";
            when "10" & x"af3" => data <= x"09";
            when "10" & x"af4" => data <= x"0d";
            when "10" & x"af5" => data <= x"a9";
            when "10" & x"af6" => data <= x"ff";
            when "10" & x"af7" => data <= x"8d";
            when "10" & x"af8" => data <= x"0a";
            when "10" & x"af9" => data <= x"0d";
            when "10" & x"afa" => data <= x"8d";
            when "10" & x"afb" => data <= x"0b";
            when "10" & x"afc" => data <= x"0d";
            when "10" & x"afd" => data <= x"4c";
            when "10" & x"afe" => data <= x"e0";
            when "10" & x"aff" => data <= x"ac";
            when "10" & x"b00" => data <= x"ad";
            when "10" & x"b01" => data <= x"fe";
            when "10" & x"b02" => data <= x"0f";
            when "10" & x"b03" => data <= x"c9";
            when "10" & x"b04" => data <= x"55";
            when "10" & x"b05" => data <= x"d0";
            when "10" & x"b06" => data <= x"05";
            when "10" & x"b07" => data <= x"ad";
            when "10" & x"b08" => data <= x"ff";
            when "10" & x"b09" => data <= x"0f";
            when "10" & x"b0a" => data <= x"c9";
            when "10" & x"b0b" => data <= x"aa";
            when "10" & x"b0c" => data <= x"60";
            when "10" & x"b0d" => data <= x"4c";
            when "10" & x"b0e" => data <= x"f1";
            when "10" & x"b0f" => data <= x"ac";
            when "10" & x"b10" => data <= x"ad";
            when "10" & x"b11" => data <= x"00";
            when "10" & x"b12" => data <= x"0e";
            when "10" & x"b13" => data <= x"c9";
            when "10" & x"b14" => data <= x"eb";
            when "10" & x"b15" => data <= x"d0";
            when "10" & x"b16" => data <= x"0e";
            when "10" & x"b17" => data <= x"ad";
            when "10" & x"b18" => data <= x"02";
            when "10" & x"b19" => data <= x"0e";
            when "10" & x"b1a" => data <= x"c9";
            when "10" & x"b1b" => data <= x"90";
            when "10" & x"b1c" => data <= x"d0";
            when "10" & x"b1d" => data <= x"07";
            when "10" & x"b1e" => data <= x"ad";
            when "10" & x"b1f" => data <= x"0c";
            when "10" & x"b20" => data <= x"0e";
            when "10" & x"b21" => data <= x"c9";
            when "10" & x"b22" => data <= x"02";
            when "10" & x"b23" => data <= x"f0";
            when "10" & x"b24" => data <= x"26";
            when "10" & x"b25" => data <= x"ad";
            when "10" & x"b26" => data <= x"c6";
            when "10" & x"b27" => data <= x"0f";
            when "10" & x"b28" => data <= x"8d";
            when "10" & x"b29" => data <= x"23";
            when "10" & x"b2a" => data <= x"0d";
            when "10" & x"b2b" => data <= x"ad";
            when "10" & x"b2c" => data <= x"c7";
            when "10" & x"b2d" => data <= x"0f";
            when "10" & x"b2e" => data <= x"8d";
            when "10" & x"b2f" => data <= x"24";
            when "10" & x"b30" => data <= x"0d";
            when "10" & x"b31" => data <= x"ad";
            when "10" & x"b32" => data <= x"c8";
            when "10" & x"b33" => data <= x"0f";
            when "10" & x"b34" => data <= x"8d";
            when "10" & x"b35" => data <= x"25";
            when "10" & x"b36" => data <= x"0d";
            when "10" & x"b37" => data <= x"ad";
            when "10" & x"b38" => data <= x"c9";
            when "10" & x"b39" => data <= x"0f";
            when "10" & x"b3a" => data <= x"8d";
            when "10" & x"b3b" => data <= x"26";
            when "10" & x"b3c" => data <= x"0d";
            when "10" & x"b3d" => data <= x"20";
            when "10" & x"b3e" => data <= x"0a";
            when "10" & x"b3f" => data <= x"ad";
            when "10" & x"b40" => data <= x"20";
            when "10" & x"b41" => data <= x"99";
            when "10" & x"b42" => data <= x"a7";
            when "10" & x"b43" => data <= x"20";
            when "10" & x"b44" => data <= x"23";
            when "10" & x"b45" => data <= x"ad";
            when "10" & x"b46" => data <= x"20";
            when "10" & x"b47" => data <= x"00";
            when "10" & x"b48" => data <= x"ab";
            when "10" & x"b49" => data <= x"d0";
            when "10" & x"b4a" => data <= x"c2";
            when "10" & x"b4b" => data <= x"ad";
            when "10" & x"b4c" => data <= x"0b";
            when "10" & x"b4d" => data <= x"0e";
            when "10" & x"b4e" => data <= x"d0";
            when "10" & x"b4f" => data <= x"bd";
            when "10" & x"b50" => data <= x"ad";
            when "10" & x"b51" => data <= x"0c";
            when "10" & x"b52" => data <= x"0e";
            when "10" & x"b53" => data <= x"c9";
            when "10" & x"b54" => data <= x"02";
            when "10" & x"b55" => data <= x"d0";
            when "10" & x"b56" => data <= x"b6";
            when "10" & x"b57" => data <= x"a2";
            when "10" & x"b58" => data <= x"05";
            when "10" & x"b59" => data <= x"0e";
            when "10" & x"b5a" => data <= x"11";
            when "10" & x"b5b" => data <= x"0e";
            when "10" & x"b5c" => data <= x"2e";
            when "10" & x"b5d" => data <= x"12";
            when "10" & x"b5e" => data <= x"0e";
            when "10" & x"b5f" => data <= x"ca";
            when "10" & x"b60" => data <= x"d0";
            when "10" & x"b61" => data <= x"f7";
            when "10" & x"b62" => data <= x"4e";
            when "10" & x"b63" => data <= x"12";
            when "10" & x"b64" => data <= x"0e";
            when "10" & x"b65" => data <= x"ad";
            when "10" & x"b66" => data <= x"12";
            when "10" & x"b67" => data <= x"0e";
            when "10" & x"b68" => data <= x"8d";
            when "10" & x"b69" => data <= x"39";
            when "10" & x"b6a" => data <= x"0d";
            when "10" & x"b6b" => data <= x"ad";
            when "10" & x"b6c" => data <= x"0d";
            when "10" & x"b6d" => data <= x"0e";
            when "10" & x"b6e" => data <= x"8d";
            when "10" & x"b6f" => data <= x"29";
            when "10" & x"b70" => data <= x"0d";
            when "10" & x"b71" => data <= x"18";
            when "10" & x"b72" => data <= x"ad";
            when "10" & x"b73" => data <= x"0e";
            when "10" & x"b74" => data <= x"0e";
            when "10" & x"b75" => data <= x"6d";
            when "10" & x"b76" => data <= x"23";
            when "10" & x"b77" => data <= x"0d";
            when "10" & x"b78" => data <= x"8d";
            when "10" & x"b79" => data <= x"23";
            when "10" & x"b7a" => data <= x"0d";
            when "10" & x"b7b" => data <= x"ad";
            when "10" & x"b7c" => data <= x"0f";
            when "10" & x"b7d" => data <= x"0e";
            when "10" & x"b7e" => data <= x"6d";
            when "10" & x"b7f" => data <= x"24";
            when "10" & x"b80" => data <= x"0d";
            when "10" & x"b81" => data <= x"8d";
            when "10" & x"b82" => data <= x"24";
            when "10" & x"b83" => data <= x"0d";
            when "10" & x"b84" => data <= x"a9";
            when "10" & x"b85" => data <= x"00";
            when "10" & x"b86" => data <= x"6d";
            when "10" & x"b87" => data <= x"25";
            when "10" & x"b88" => data <= x"0d";
            when "10" & x"b89" => data <= x"8d";
            when "10" & x"b8a" => data <= x"25";
            when "10" & x"b8b" => data <= x"0d";
            when "10" & x"b8c" => data <= x"a9";
            when "10" & x"b8d" => data <= x"00";
            when "10" & x"b8e" => data <= x"6d";
            when "10" & x"b8f" => data <= x"26";
            when "10" & x"b90" => data <= x"0d";
            when "10" & x"b91" => data <= x"8d";
            when "10" & x"b92" => data <= x"26";
            when "10" & x"b93" => data <= x"0d";
            when "10" & x"b94" => data <= x"90";
            when "10" & x"b95" => data <= x"03";
            when "10" & x"b96" => data <= x"4c";
            when "10" & x"b97" => data <= x"f1";
            when "10" & x"b98" => data <= x"ac";
            when "10" & x"b99" => data <= x"ad";
            when "10" & x"b9a" => data <= x"11";
            when "10" & x"b9b" => data <= x"0e";
            when "10" & x"b9c" => data <= x"0d";
            when "10" & x"b9d" => data <= x"12";
            when "10" & x"b9e" => data <= x"0e";
            when "10" & x"b9f" => data <= x"8d";
            when "10" & x"ba0" => data <= x"22";
            when "10" & x"ba1" => data <= x"0d";
            when "10" & x"ba2" => data <= x"f0";
            when "10" & x"ba3" => data <= x"14";
            when "10" & x"ba4" => data <= x"a9";
            when "10" & x"ba5" => data <= x"00";
            when "10" & x"ba6" => data <= x"8d";
            when "10" & x"ba7" => data <= x"26";
            when "10" & x"ba8" => data <= x"0e";
            when "10" & x"ba9" => data <= x"8d";
            when "10" & x"baa" => data <= x"27";
            when "10" & x"bab" => data <= x"0e";
            when "10" & x"bac" => data <= x"ad";
            when "10" & x"bad" => data <= x"16";
            when "10" & x"bae" => data <= x"0e";
            when "10" & x"baf" => data <= x"8d";
            when "10" & x"bb0" => data <= x"24";
            when "10" & x"bb1" => data <= x"0e";
            when "10" & x"bb2" => data <= x"ad";
            when "10" & x"bb3" => data <= x"17";
            when "10" & x"bb4" => data <= x"0e";
            when "10" & x"bb5" => data <= x"8d";
            when "10" & x"bb6" => data <= x"25";
            when "10" & x"bb7" => data <= x"0e";
            when "10" & x"bb8" => data <= x"ae";
            when "10" & x"bb9" => data <= x"10";
            when "10" & x"bba" => data <= x"0e";
            when "10" & x"bbb" => data <= x"18";
            when "10" & x"bbc" => data <= x"ad";
            when "10" & x"bbd" => data <= x"23";
            when "10" & x"bbe" => data <= x"0d";
            when "10" & x"bbf" => data <= x"6d";
            when "10" & x"bc0" => data <= x"24";
            when "10" & x"bc1" => data <= x"0e";
            when "10" & x"bc2" => data <= x"8d";
            when "10" & x"bc3" => data <= x"23";
            when "10" & x"bc4" => data <= x"0d";
            when "10" & x"bc5" => data <= x"ad";
            when "10" & x"bc6" => data <= x"24";
            when "10" & x"bc7" => data <= x"0d";
            when "10" & x"bc8" => data <= x"6d";
            when "10" & x"bc9" => data <= x"25";
            when "10" & x"bca" => data <= x"0e";
            when "10" & x"bcb" => data <= x"8d";
            when "10" & x"bcc" => data <= x"24";
            when "10" & x"bcd" => data <= x"0d";
            when "10" & x"bce" => data <= x"ad";
            when "10" & x"bcf" => data <= x"25";
            when "10" & x"bd0" => data <= x"0d";
            when "10" & x"bd1" => data <= x"6d";
            when "10" & x"bd2" => data <= x"26";
            when "10" & x"bd3" => data <= x"0e";
            when "10" & x"bd4" => data <= x"8d";
            when "10" & x"bd5" => data <= x"25";
            when "10" & x"bd6" => data <= x"0d";
            when "10" & x"bd7" => data <= x"ad";
            when "10" & x"bd8" => data <= x"26";
            when "10" & x"bd9" => data <= x"0d";
            when "10" & x"bda" => data <= x"6d";
            when "10" & x"bdb" => data <= x"27";
            when "10" & x"bdc" => data <= x"0e";
            when "10" & x"bdd" => data <= x"8d";
            when "10" & x"bde" => data <= x"26";
            when "10" & x"bdf" => data <= x"0d";
            when "10" & x"be0" => data <= x"90";
            when "10" & x"be1" => data <= x"03";
            when "10" & x"be2" => data <= x"4c";
            when "10" & x"be3" => data <= x"0d";
            when "10" & x"be4" => data <= x"ab";
            when "10" & x"be5" => data <= x"ca";
            when "10" & x"be6" => data <= x"d0";
            when "10" & x"be7" => data <= x"d3";
            when "10" & x"be8" => data <= x"a9";
            when "10" & x"be9" => data <= x"20";
            when "10" & x"bea" => data <= x"8d";
            when "10" & x"beb" => data <= x"21";
            when "10" & x"bec" => data <= x"0d";
            when "10" & x"bed" => data <= x"20";
            when "10" & x"bee" => data <= x"0a";
            when "10" & x"bef" => data <= x"ad";
            when "10" & x"bf0" => data <= x"20";
            when "10" & x"bf1" => data <= x"99";
            when "10" & x"bf2" => data <= x"a7";
            when "10" & x"bf3" => data <= x"20";
            when "10" & x"bf4" => data <= x"23";
            when "10" & x"bf5" => data <= x"ad";
            when "10" & x"bf6" => data <= x"a9";
            when "10" & x"bf7" => data <= x"00";
            when "10" & x"bf8" => data <= x"85";
            when "10" & x"bf9" => data <= x"a2";
            when "10" & x"bfa" => data <= x"a9";
            when "10" & x"bfb" => data <= x"0e";
            when "10" & x"bfc" => data <= x"85";
            when "10" & x"bfd" => data <= x"a3";
            when "10" & x"bfe" => data <= x"a0";
            when "10" & x"bff" => data <= x"0b";
            when "10" & x"c00" => data <= x"b1";
            when "10" & x"c01" => data <= x"a2";
            when "10" & x"c02" => data <= x"29";
            when "10" & x"c03" => data <= x"0f";
            when "10" & x"c04" => data <= x"d0";
            when "10" & x"c05" => data <= x"10";
            when "10" & x"c06" => data <= x"a0";
            when "10" & x"c07" => data <= x"00";
            when "10" & x"c08" => data <= x"b1";
            when "10" & x"c09" => data <= x"a2";
            when "10" & x"c0a" => data <= x"d9";
            when "10" & x"c0b" => data <= x"70";
            when "10" & x"c0c" => data <= x"0d";
            when "10" & x"c0d" => data <= x"d0";
            when "10" & x"c0e" => data <= x"07";
            when "10" & x"c0f" => data <= x"c8";
            when "10" & x"c10" => data <= x"c0";
            when "10" & x"c11" => data <= x"0b";
            when "10" & x"c12" => data <= x"f0";
            when "10" & x"c13" => data <= x"38";
            when "10" & x"c14" => data <= x"d0";
            when "10" & x"c15" => data <= x"f2";
            when "10" & x"c16" => data <= x"18";
            when "10" & x"c17" => data <= x"a5";
            when "10" & x"c18" => data <= x"a2";
            when "10" & x"c19" => data <= x"69";
            when "10" & x"c1a" => data <= x"20";
            when "10" & x"c1b" => data <= x"85";
            when "10" & x"c1c" => data <= x"a2";
            when "10" & x"c1d" => data <= x"d0";
            when "10" & x"c1e" => data <= x"df";
            when "10" & x"c1f" => data <= x"e6";
            when "10" & x"c20" => data <= x"a3";
            when "10" & x"c21" => data <= x"a5";
            when "10" & x"c22" => data <= x"a3";
            when "10" & x"c23" => data <= x"c9";
            when "10" & x"c24" => data <= x"0f";
            when "10" & x"c25" => data <= x"f0";
            when "10" & x"c26" => data <= x"d7";
            when "10" & x"c27" => data <= x"ce";
            when "10" & x"c28" => data <= x"21";
            when "10" & x"c29" => data <= x"0d";
            when "10" & x"c2a" => data <= x"ad";
            when "10" & x"c2b" => data <= x"21";
            when "10" & x"c2c" => data <= x"0d";
            when "10" & x"c2d" => data <= x"f0";
            when "10" & x"c2e" => data <= x"08";
            when "10" & x"c2f" => data <= x"a9";
            when "10" & x"c30" => data <= x"01";
            when "10" & x"c31" => data <= x"20";
            when "10" & x"c32" => data <= x"3c";
            when "10" & x"c33" => data <= x"ad";
            when "10" & x"c34" => data <= x"4c";
            when "10" & x"c35" => data <= x"ed";
            when "10" & x"c36" => data <= x"ab";
            when "10" & x"c37" => data <= x"20";
            when "10" & x"c38" => data <= x"00";
            when "10" & x"c39" => data <= x"a0";
            when "10" & x"c3a" => data <= x"ff";
            when "10" & x"c3b" => data <= x"49";
            when "10" & x"c3c" => data <= x"6d";
            when "10" & x"c3d" => data <= x"61";
            when "10" & x"c3e" => data <= x"67";
            when "10" & x"c3f" => data <= x"65";
            when "10" & x"c40" => data <= x"20";
            when "10" & x"c41" => data <= x"6e";
            when "10" & x"c42" => data <= x"6f";
            when "10" & x"c43" => data <= x"74";
            when "10" & x"c44" => data <= x"20";
            when "10" & x"c45" => data <= x"66";
            when "10" & x"c46" => data <= x"6f";
            when "10" & x"c47" => data <= x"75";
            when "10" & x"c48" => data <= x"6e";
            when "10" & x"c49" => data <= x"64";
            when "10" & x"c4a" => data <= x"21";
            when "10" & x"c4b" => data <= x"00";
            when "10" & x"c4c" => data <= x"a0";
            when "10" & x"c4d" => data <= x"14";
            when "10" & x"c4e" => data <= x"b1";
            when "10" & x"c4f" => data <= x"a2";
            when "10" & x"c50" => data <= x"8d";
            when "10" & x"c51" => data <= x"2c";
            when "10" & x"c52" => data <= x"0d";
            when "10" & x"c53" => data <= x"c8";
            when "10" & x"c54" => data <= x"b1";
            when "10" & x"c55" => data <= x"a2";
            when "10" & x"c56" => data <= x"8d";
            when "10" & x"c57" => data <= x"2d";
            when "10" & x"c58" => data <= x"0d";
            when "10" & x"c59" => data <= x"a0";
            when "10" & x"c5a" => data <= x"1b";
            when "10" & x"c5b" => data <= x"b1";
            when "10" & x"c5c" => data <= x"a2";
            when "10" & x"c5d" => data <= x"48";
            when "10" & x"c5e" => data <= x"88";
            when "10" & x"c5f" => data <= x"b1";
            when "10" & x"c60" => data <= x"a2";
            when "10" & x"c61" => data <= x"38";
            when "10" & x"c62" => data <= x"e9";
            when "10" & x"c63" => data <= x"02";
            when "10" & x"c64" => data <= x"8d";
            when "10" & x"c65" => data <= x"2a";
            when "10" & x"c66" => data <= x"0d";
            when "10" & x"c67" => data <= x"68";
            when "10" & x"c68" => data <= x"e9";
            when "10" & x"c69" => data <= x"00";
            when "10" & x"c6a" => data <= x"8d";
            when "10" & x"c6b" => data <= x"2b";
            when "10" & x"c6c" => data <= x"0d";
            when "10" & x"c6d" => data <= x"ad";
            when "10" & x"c6e" => data <= x"2c";
            when "10" & x"c6f" => data <= x"0d";
            when "10" & x"c70" => data <= x"e9";
            when "10" & x"c71" => data <= x"00";
            when "10" & x"c72" => data <= x"8d";
            when "10" & x"c73" => data <= x"2c";
            when "10" & x"c74" => data <= x"0d";
            when "10" & x"c75" => data <= x"ad";
            when "10" & x"c76" => data <= x"2d";
            when "10" & x"c77" => data <= x"0d";
            when "10" & x"c78" => data <= x"e9";
            when "10" & x"c79" => data <= x"00";
            when "10" & x"c7a" => data <= x"8d";
            when "10" & x"c7b" => data <= x"2d";
            when "10" & x"c7c" => data <= x"0d";
            when "10" & x"c7d" => data <= x"0d";
            when "10" & x"c7e" => data <= x"2c";
            when "10" & x"c7f" => data <= x"0d";
            when "10" & x"c80" => data <= x"0d";
            when "10" & x"c81" => data <= x"2b";
            when "10" & x"c82" => data <= x"0d";
            when "10" & x"c83" => data <= x"0d";
            when "10" & x"c84" => data <= x"2a";
            when "10" & x"c85" => data <= x"0d";
            when "10" & x"c86" => data <= x"f0";
            when "10" & x"c87" => data <= x"2b";
            when "10" & x"c88" => data <= x"ae";
            when "10" & x"c89" => data <= x"29";
            when "10" & x"c8a" => data <= x"0d";
            when "10" & x"c8b" => data <= x"18";
            when "10" & x"c8c" => data <= x"ad";
            when "10" & x"c8d" => data <= x"23";
            when "10" & x"c8e" => data <= x"0d";
            when "10" & x"c8f" => data <= x"6d";
            when "10" & x"c90" => data <= x"2a";
            when "10" & x"c91" => data <= x"0d";
            when "10" & x"c92" => data <= x"8d";
            when "10" & x"c93" => data <= x"23";
            when "10" & x"c94" => data <= x"0d";
            when "10" & x"c95" => data <= x"ad";
            when "10" & x"c96" => data <= x"24";
            when "10" & x"c97" => data <= x"0d";
            when "10" & x"c98" => data <= x"6d";
            when "10" & x"c99" => data <= x"2b";
            when "10" & x"c9a" => data <= x"0d";
            when "10" & x"c9b" => data <= x"8d";
            when "10" & x"c9c" => data <= x"24";
            when "10" & x"c9d" => data <= x"0d";
            when "10" & x"c9e" => data <= x"ad";
            when "10" & x"c9f" => data <= x"25";
            when "10" & x"ca0" => data <= x"0d";
            when "10" & x"ca1" => data <= x"6d";
            when "10" & x"ca2" => data <= x"2c";
            when "10" & x"ca3" => data <= x"0d";
            when "10" & x"ca4" => data <= x"8d";
            when "10" & x"ca5" => data <= x"25";
            when "10" & x"ca6" => data <= x"0d";
            when "10" & x"ca7" => data <= x"ad";
            when "10" & x"ca8" => data <= x"26";
            when "10" & x"ca9" => data <= x"0d";
            when "10" & x"caa" => data <= x"6d";
            when "10" & x"cab" => data <= x"2d";
            when "10" & x"cac" => data <= x"0d";
            when "10" & x"cad" => data <= x"8d";
            when "10" & x"cae" => data <= x"26";
            when "10" & x"caf" => data <= x"0d";
            when "10" & x"cb0" => data <= x"ca";
            when "10" & x"cb1" => data <= x"d0";
            when "10" & x"cb2" => data <= x"d8";
            when "10" & x"cb3" => data <= x"ad";
            when "10" & x"cb4" => data <= x"22";
            when "10" & x"cb5" => data <= x"0d";
            when "10" & x"cb6" => data <= x"f0";
            when "10" & x"cb7" => data <= x"06";
            when "10" & x"cb8" => data <= x"ad";
            when "10" & x"cb9" => data <= x"39";
            when "10" & x"cba" => data <= x"0d";
            when "10" & x"cbb" => data <= x"20";
            when "10" & x"cbc" => data <= x"3c";
            when "10" & x"cbd" => data <= x"ad";
            when "10" & x"cbe" => data <= x"ad";
            when "10" & x"cbf" => data <= x"23";
            when "10" & x"cc0" => data <= x"0d";
            when "10" & x"cc1" => data <= x"8d";
            when "10" & x"cc2" => data <= x"06";
            when "10" & x"cc3" => data <= x"0d";
            when "10" & x"cc4" => data <= x"49";
            when "10" & x"cc5" => data <= x"ff";
            when "10" & x"cc6" => data <= x"8d";
            when "10" & x"cc7" => data <= x"0a";
            when "10" & x"cc8" => data <= x"0d";
            when "10" & x"cc9" => data <= x"ad";
            when "10" & x"cca" => data <= x"24";
            when "10" & x"ccb" => data <= x"0d";
            when "10" & x"ccc" => data <= x"8d";
            when "10" & x"ccd" => data <= x"07";
            when "10" & x"cce" => data <= x"0d";
            when "10" & x"ccf" => data <= x"49";
            when "10" & x"cd0" => data <= x"ff";
            when "10" & x"cd1" => data <= x"8d";
            when "10" & x"cd2" => data <= x"0b";
            when "10" & x"cd3" => data <= x"0d";
            when "10" & x"cd4" => data <= x"ad";
            when "10" & x"cd5" => data <= x"25";
            when "10" & x"cd6" => data <= x"0d";
            when "10" & x"cd7" => data <= x"8d";
            when "10" & x"cd8" => data <= x"08";
            when "10" & x"cd9" => data <= x"0d";
            when "10" & x"cda" => data <= x"ad";
            when "10" & x"cdb" => data <= x"26";
            when "10" & x"cdc" => data <= x"0d";
            when "10" & x"cdd" => data <= x"8d";
            when "10" & x"cde" => data <= x"09";
            when "10" & x"cdf" => data <= x"0d";
            when "10" & x"ce0" => data <= x"a9";
            when "10" & x"ce1" => data <= x"54";
            when "10" & x"ce2" => data <= x"8d";
            when "10" & x"ce3" => data <= x"05";
            when "10" & x"ce4" => data <= x"0d";
            when "10" & x"ce5" => data <= x"a2";
            when "10" & x"ce6" => data <= x"00";
            when "10" & x"ce7" => data <= x"68";
            when "10" & x"ce8" => data <= x"9d";
            when "10" & x"ce9" => data <= x"23";
            when "10" & x"cea" => data <= x"0d";
            when "10" & x"ceb" => data <= x"e8";
            when "10" & x"cec" => data <= x"e0";
            when "10" & x"ced" => data <= x"0b";
            when "10" & x"cee" => data <= x"d0";
            when "10" & x"cef" => data <= x"f7";
            when "10" & x"cf0" => data <= x"60";
            when "10" & x"cf1" => data <= x"20";
            when "10" & x"cf2" => data <= x"00";
            when "10" & x"cf3" => data <= x"a0";
            when "10" & x"cf4" => data <= x"ff";
            when "10" & x"cf5" => data <= x"55";
            when "10" & x"cf6" => data <= x"6e";
            when "10" & x"cf7" => data <= x"72";
            when "10" & x"cf8" => data <= x"65";
            when "10" & x"cf9" => data <= x"63";
            when "10" & x"cfa" => data <= x"6f";
            when "10" & x"cfb" => data <= x"67";
            when "10" & x"cfc" => data <= x"6e";
            when "10" & x"cfd" => data <= x"69";
            when "10" & x"cfe" => data <= x"73";
            when "10" & x"cff" => data <= x"65";
            when "10" & x"d00" => data <= x"64";
            when "10" & x"d01" => data <= x"20";
            when "10" & x"d02" => data <= x"66";
            when "10" & x"d03" => data <= x"6f";
            when "10" & x"d04" => data <= x"72";
            when "10" & x"d05" => data <= x"6d";
            when "10" & x"d06" => data <= x"61";
            when "10" & x"d07" => data <= x"74";
            when "10" & x"d08" => data <= x"21";
            when "10" & x"d09" => data <= x"00";
            when "10" & x"d0a" => data <= x"ad";
            when "10" & x"d0b" => data <= x"23";
            when "10" & x"d0c" => data <= x"0d";
            when "10" & x"d0d" => data <= x"8d";
            when "10" & x"d0e" => data <= x"06";
            when "10" & x"d0f" => data <= x"0d";
            when "10" & x"d10" => data <= x"ad";
            when "10" & x"d11" => data <= x"24";
            when "10" & x"d12" => data <= x"0d";
            when "10" & x"d13" => data <= x"8d";
            when "10" & x"d14" => data <= x"07";
            when "10" & x"d15" => data <= x"0d";
            when "10" & x"d16" => data <= x"ad";
            when "10" & x"d17" => data <= x"25";
            when "10" & x"d18" => data <= x"0d";
            when "10" & x"d19" => data <= x"8d";
            when "10" & x"d1a" => data <= x"08";
            when "10" & x"d1b" => data <= x"0d";
            when "10" & x"d1c" => data <= x"ad";
            when "10" & x"d1d" => data <= x"26";
            when "10" & x"d1e" => data <= x"0d";
            when "10" & x"d1f" => data <= x"8d";
            when "10" & x"d20" => data <= x"09";
            when "10" & x"d21" => data <= x"0d";
            when "10" & x"d22" => data <= x"60";
            when "10" & x"d23" => data <= x"ad";
            when "10" & x"d24" => data <= x"06";
            when "10" & x"d25" => data <= x"0d";
            when "10" & x"d26" => data <= x"8d";
            when "10" & x"d27" => data <= x"23";
            when "10" & x"d28" => data <= x"0d";
            when "10" & x"d29" => data <= x"ad";
            when "10" & x"d2a" => data <= x"07";
            when "10" & x"d2b" => data <= x"0d";
            when "10" & x"d2c" => data <= x"8d";
            when "10" & x"d2d" => data <= x"24";
            when "10" & x"d2e" => data <= x"0d";
            when "10" & x"d2f" => data <= x"ad";
            when "10" & x"d30" => data <= x"08";
            when "10" & x"d31" => data <= x"0d";
            when "10" & x"d32" => data <= x"8d";
            when "10" & x"d33" => data <= x"25";
            when "10" & x"d34" => data <= x"0d";
            when "10" & x"d35" => data <= x"ad";
            when "10" & x"d36" => data <= x"09";
            when "10" & x"d37" => data <= x"0d";
            when "10" & x"d38" => data <= x"8d";
            when "10" & x"d39" => data <= x"26";
            when "10" & x"d3a" => data <= x"0d";
            when "10" & x"d3b" => data <= x"60";
            when "10" & x"d3c" => data <= x"18";
            when "10" & x"d3d" => data <= x"6d";
            when "10" & x"d3e" => data <= x"23";
            when "10" & x"d3f" => data <= x"0d";
            when "10" & x"d40" => data <= x"8d";
            when "10" & x"d41" => data <= x"23";
            when "10" & x"d42" => data <= x"0d";
            when "10" & x"d43" => data <= x"ad";
            when "10" & x"d44" => data <= x"24";
            when "10" & x"d45" => data <= x"0d";
            when "10" & x"d46" => data <= x"69";
            when "10" & x"d47" => data <= x"00";
            when "10" & x"d48" => data <= x"8d";
            when "10" & x"d49" => data <= x"24";
            when "10" & x"d4a" => data <= x"0d";
            when "10" & x"d4b" => data <= x"ad";
            when "10" & x"d4c" => data <= x"25";
            when "10" & x"d4d" => data <= x"0d";
            when "10" & x"d4e" => data <= x"69";
            when "10" & x"d4f" => data <= x"00";
            when "10" & x"d50" => data <= x"8d";
            when "10" & x"d51" => data <= x"25";
            when "10" & x"d52" => data <= x"0d";
            when "10" & x"d53" => data <= x"ad";
            when "10" & x"d54" => data <= x"26";
            when "10" & x"d55" => data <= x"0d";
            when "10" & x"d56" => data <= x"69";
            when "10" & x"d57" => data <= x"00";
            when "10" & x"d58" => data <= x"8d";
            when "10" & x"d59" => data <= x"26";
            when "10" & x"d5a" => data <= x"0d";
            when "10" & x"d5b" => data <= x"90";
            when "10" & x"d5c" => data <= x"03";
            when "10" & x"d5d" => data <= x"4c";
            when "10" & x"d5e" => data <= x"f1";
            when "10" & x"d5f" => data <= x"ac";
            when "10" & x"d60" => data <= x"60";
            when "10" & x"d61" => data <= x"42";
            when "10" & x"d62" => data <= x"45";
            when "10" & x"d63" => data <= x"45";
            when "10" & x"d64" => data <= x"42";
            when "10" & x"d65" => data <= x"20";
            when "10" & x"d66" => data <= x"20";
            when "10" & x"d67" => data <= x"20";
            when "10" & x"d68" => data <= x"20";
            when "10" & x"d69" => data <= x"4d";
            when "10" & x"d6a" => data <= x"4d";
            when "10" & x"d6b" => data <= x"42";
            when "10" & x"d6c" => data <= x"08";
            when "10" & x"d6d" => data <= x"aa";
            when "10" & x"d6e" => data <= x"20";
            when "10" & x"d6f" => data <= x"a1";
            when "10" & x"d70" => data <= x"ad";
            when "10" & x"d71" => data <= x"85";
            when "10" & x"d72" => data <= x"b2";
            when "10" & x"d73" => data <= x"48";
            when "10" & x"d74" => data <= x"20";
            when "10" & x"d75" => data <= x"bd";
            when "10" & x"d76" => data <= x"ad";
            when "10" & x"d77" => data <= x"8a";
            when "10" & x"d78" => data <= x"e5";
            when "10" & x"d79" => data <= x"b0";
            when "10" & x"d7a" => data <= x"aa";
            when "10" & x"d7b" => data <= x"68";
            when "10" & x"d7c" => data <= x"20";
            when "10" & x"d7d" => data <= x"a1";
            when "10" & x"d7e" => data <= x"ad";
            when "10" & x"d7f" => data <= x"48";
            when "10" & x"d80" => data <= x"20";
            when "10" & x"d81" => data <= x"bd";
            when "10" & x"d82" => data <= x"ad";
            when "10" & x"d83" => data <= x"a5";
            when "10" & x"d84" => data <= x"b2";
            when "10" & x"d85" => data <= x"e5";
            when "10" & x"d86" => data <= x"b0";
            when "10" & x"d87" => data <= x"0a";
            when "10" & x"d88" => data <= x"0a";
            when "10" & x"d89" => data <= x"0a";
            when "10" & x"d8a" => data <= x"0a";
            when "10" & x"d8b" => data <= x"85";
            when "10" & x"d8c" => data <= x"b2";
            when "10" & x"d8d" => data <= x"8a";
            when "10" & x"d8e" => data <= x"05";
            when "10" & x"d8f" => data <= x"b2";
            when "10" & x"d90" => data <= x"aa";
            when "10" & x"d91" => data <= x"68";
            when "10" & x"d92" => data <= x"28";
            when "10" & x"d93" => data <= x"90";
            when "10" & x"d94" => data <= x"0b";
            when "10" & x"d95" => data <= x"48";
            when "10" & x"d96" => data <= x"8a";
            when "10" & x"d97" => data <= x"f8";
            when "10" & x"d98" => data <= x"18";
            when "10" & x"d99" => data <= x"69";
            when "10" & x"d9a" => data <= x"56";
            when "10" & x"d9b" => data <= x"aa";
            when "10" & x"d9c" => data <= x"68";
            when "10" & x"d9d" => data <= x"69";
            when "10" & x"d9e" => data <= x"02";
            when "10" & x"d9f" => data <= x"d8";
            when "10" & x"da0" => data <= x"60";
            when "10" & x"da1" => data <= x"a0";
            when "10" & x"da2" => data <= x"00";
            when "10" & x"da3" => data <= x"84";
            when "10" & x"da4" => data <= x"b1";
            when "10" & x"da5" => data <= x"a0";
            when "10" & x"da6" => data <= x"a0";
            when "10" & x"da7" => data <= x"84";
            when "10" & x"da8" => data <= x"b0";
            when "10" & x"da9" => data <= x"a0";
            when "10" & x"daa" => data <= x"05";
            when "10" & x"dab" => data <= x"c5";
            when "10" & x"dac" => data <= x"b0";
            when "10" & x"dad" => data <= x"90";
            when "10" & x"dae" => data <= x"04";
            when "10" & x"daf" => data <= x"38";
            when "10" & x"db0" => data <= x"e5";
            when "10" & x"db1" => data <= x"b0";
            when "10" & x"db2" => data <= x"38";
            when "10" & x"db3" => data <= x"26";
            when "10" & x"db4" => data <= x"b1";
            when "10" & x"db5" => data <= x"46";
            when "10" & x"db6" => data <= x"b0";
            when "10" & x"db7" => data <= x"88";
            when "10" & x"db8" => data <= x"d0";
            when "10" & x"db9" => data <= x"f1";
            when "10" & x"dba" => data <= x"a5";
            when "10" & x"dbb" => data <= x"b1";
            when "10" & x"dbc" => data <= x"60";
            when "10" & x"dbd" => data <= x"48";
            when "10" & x"dbe" => data <= x"0a";
            when "10" & x"dbf" => data <= x"0a";
            when "10" & x"dc0" => data <= x"0a";
            when "10" & x"dc1" => data <= x"85";
            when "10" & x"dc2" => data <= x"b0";
            when "10" & x"dc3" => data <= x"68";
            when "10" & x"dc4" => data <= x"0a";
            when "10" & x"dc5" => data <= x"18";
            when "10" & x"dc6" => data <= x"65";
            when "10" & x"dc7" => data <= x"b0";
            when "10" & x"dc8" => data <= x"85";
            when "10" & x"dc9" => data <= x"b0";
            when "10" & x"dca" => data <= x"38";
            when "10" & x"dcb" => data <= x"60";
            when "10" & x"dcc" => data <= x"e0";
            when "10" & x"dcd" => data <= x"ff";
            when "10" & x"dce" => data <= x"f0";
            when "10" & x"dcf" => data <= x"35";
            when "10" & x"dd0" => data <= x"bd";
            when "10" & x"dd1" => data <= x"10";
            when "10" & x"dd2" => data <= x"0d";
            when "10" & x"dd3" => data <= x"30";
            when "10" & x"dd4" => data <= x"30";
            when "10" & x"dd5" => data <= x"49";
            when "10" & x"dd6" => data <= x"ff";
            when "10" & x"dd7" => data <= x"dd";
            when "10" & x"dd8" => data <= x"18";
            when "10" & x"dd9" => data <= x"0d";
            when "10" & x"dda" => data <= x"d0";
            when "10" & x"ddb" => data <= x"24";
            when "10" & x"ddc" => data <= x"bd";
            when "10" & x"ddd" => data <= x"0c";
            when "10" & x"dde" => data <= x"0d";
            when "10" & x"ddf" => data <= x"49";
            when "10" & x"de0" => data <= x"ff";
            when "10" & x"de1" => data <= x"dd";
            when "10" & x"de2" => data <= x"14";
            when "10" & x"de3" => data <= x"0d";
            when "10" & x"de4" => data <= x"d0";
            when "10" & x"de5" => data <= x"1a";
            when "10" & x"de6" => data <= x"bd";
            when "10" & x"de7" => data <= x"1c";
            when "10" & x"de8" => data <= x"0d";
            when "10" & x"de9" => data <= x"c9";
            when "10" & x"dea" => data <= x"54";
            when "10" & x"deb" => data <= x"f0";
            when "10" & x"dec" => data <= x"29";
            when "10" & x"ded" => data <= x"20";
            when "10" & x"dee" => data <= x"00";
            when "10" & x"def" => data <= x"a0";
            when "10" & x"df0" => data <= x"c9";
            when "10" & x"df1" => data <= x"44";
            when "10" & x"df2" => data <= x"69";
            when "10" & x"df3" => data <= x"73";
            when "10" & x"df4" => data <= x"6b";
            when "10" & x"df5" => data <= x"20";
            when "10" & x"df6" => data <= x"72";
            when "10" & x"df7" => data <= x"65";
            when "10" & x"df8" => data <= x"61";
            when "10" & x"df9" => data <= x"64";
            when "10" & x"dfa" => data <= x"20";
            when "10" & x"dfb" => data <= x"6f";
            when "10" & x"dfc" => data <= x"6e";
            when "10" & x"dfd" => data <= x"6c";
            when "10" & x"dfe" => data <= x"79";
            when "10" & x"dff" => data <= x"00";
            when "10" & x"e00" => data <= x"a9";
            when "10" & x"e01" => data <= x"ff";
            when "10" & x"e02" => data <= x"9d";
            when "10" & x"e03" => data <= x"10";
            when "10" & x"e04" => data <= x"0d";
            when "10" & x"e05" => data <= x"20";
            when "10" & x"e06" => data <= x"00";
            when "10" & x"e07" => data <= x"a0";
            when "10" & x"e08" => data <= x"c7";
            when "10" & x"e09" => data <= x"4e";
            when "10" & x"e0a" => data <= x"6f";
            when "10" & x"e0b" => data <= x"20";
            when "10" & x"e0c" => data <= x"64";
            when "10" & x"e0d" => data <= x"69";
            when "10" & x"e0e" => data <= x"73";
            when "10" & x"e0f" => data <= x"6b";
            when "10" & x"e10" => data <= x"00";
            when "10" & x"e11" => data <= x"a9";
            when "10" & x"e12" => data <= x"54";
            when "10" & x"e13" => data <= x"9d";
            when "10" & x"e14" => data <= x"1c";
            when "10" & x"e15" => data <= x"0d";
            when "10" & x"e16" => data <= x"60";
            when "10" & x"e17" => data <= x"a9";
            when "10" & x"e18" => data <= x"00";
            when "10" & x"e19" => data <= x"9d";
            when "10" & x"e1a" => data <= x"1c";
            when "10" & x"e1b" => data <= x"0d";
            when "10" & x"e1c" => data <= x"60";
            when "10" & x"e1d" => data <= x"bd";
            when "10" & x"e1e" => data <= x"10";
            when "10" & x"e1f" => data <= x"0d";
            when "10" & x"e20" => data <= x"30";
            when "10" & x"e21" => data <= x"e3";
            when "10" & x"e22" => data <= x"6a";
            when "10" & x"e23" => data <= x"bd";
            when "10" & x"e24" => data <= x"0c";
            when "10" & x"e25" => data <= x"0d";
            when "10" & x"e26" => data <= x"08";
            when "10" & x"e27" => data <= x"aa";
            when "10" & x"e28" => data <= x"a9";
            when "10" & x"e29" => data <= x"00";
            when "10" & x"e2a" => data <= x"8d";
            when "10" & x"e2b" => data <= x"23";
            when "10" & x"e2c" => data <= x"0d";
            when "10" & x"e2d" => data <= x"8d";
            when "10" & x"e2e" => data <= x"26";
            when "10" & x"e2f" => data <= x"0d";
            when "10" & x"e30" => data <= x"2a";
            when "10" & x"e31" => data <= x"48";
            when "10" & x"e32" => data <= x"8d";
            when "10" & x"e33" => data <= x"25";
            when "10" & x"e34" => data <= x"0d";
            when "10" & x"e35" => data <= x"8a";
            when "10" & x"e36" => data <= x"0a";
            when "10" & x"e37" => data <= x"2e";
            when "10" & x"e38" => data <= x"25";
            when "10" & x"e39" => data <= x"0d";
            when "10" & x"e3a" => data <= x"8d";
            when "10" & x"e3b" => data <= x"24";
            when "10" & x"e3c" => data <= x"0d";
            when "10" & x"e3d" => data <= x"8a";
            when "10" & x"e3e" => data <= x"6d";
            when "10" & x"e3f" => data <= x"24";
            when "10" & x"e40" => data <= x"0d";
            when "10" & x"e41" => data <= x"8d";
            when "10" & x"e42" => data <= x"24";
            when "10" & x"e43" => data <= x"0d";
            when "10" & x"e44" => data <= x"68";
            when "10" & x"e45" => data <= x"69";
            when "10" & x"e46" => data <= x"00";
            when "10" & x"e47" => data <= x"6d";
            when "10" & x"e48" => data <= x"25";
            when "10" & x"e49" => data <= x"0d";
            when "10" & x"e4a" => data <= x"8d";
            when "10" & x"e4b" => data <= x"25";
            when "10" & x"e4c" => data <= x"0d";
            when "10" & x"e4d" => data <= x"a9";
            when "10" & x"e4e" => data <= x"00";
            when "10" & x"e4f" => data <= x"6d";
            when "10" & x"e50" => data <= x"26";
            when "10" & x"e51" => data <= x"0d";
            when "10" & x"e52" => data <= x"8d";
            when "10" & x"e53" => data <= x"26";
            when "10" & x"e54" => data <= x"0d";
            when "10" & x"e55" => data <= x"6e";
            when "10" & x"e56" => data <= x"23";
            when "10" & x"e57" => data <= x"0d";
            when "10" & x"e58" => data <= x"8a";
            when "10" & x"e59" => data <= x"28";
            when "10" & x"e5a" => data <= x"6a";
            when "10" & x"e5b" => data <= x"6e";
            when "10" & x"e5c" => data <= x"23";
            when "10" & x"e5d" => data <= x"0d";
            when "10" & x"e5e" => data <= x"4a";
            when "10" & x"e5f" => data <= x"6e";
            when "10" & x"e60" => data <= x"23";
            when "10" & x"e61" => data <= x"0d";
            when "10" & x"e62" => data <= x"4a";
            when "10" & x"e63" => data <= x"6e";
            when "10" & x"e64" => data <= x"23";
            when "10" & x"e65" => data <= x"0d";
            when "10" & x"e66" => data <= x"6d";
            when "10" & x"e67" => data <= x"24";
            when "10" & x"e68" => data <= x"0d";
            when "10" & x"e69" => data <= x"8d";
            when "10" & x"e6a" => data <= x"24";
            when "10" & x"e6b" => data <= x"0d";
            when "10" & x"e6c" => data <= x"ad";
            when "10" & x"e6d" => data <= x"25";
            when "10" & x"e6e" => data <= x"0d";
            when "10" & x"e6f" => data <= x"69";
            when "10" & x"e70" => data <= x"00";
            when "10" & x"e71" => data <= x"8d";
            when "10" & x"e72" => data <= x"25";
            when "10" & x"e73" => data <= x"0d";
            when "10" & x"e74" => data <= x"ad";
            when "10" & x"e75" => data <= x"26";
            when "10" & x"e76" => data <= x"0d";
            when "10" & x"e77" => data <= x"69";
            when "10" & x"e78" => data <= x"00";
            when "10" & x"e79" => data <= x"8d";
            when "10" & x"e7a" => data <= x"26";
            when "10" & x"e7b" => data <= x"0d";
            when "10" & x"e7c" => data <= x"6e";
            when "10" & x"e7d" => data <= x"26";
            when "10" & x"e7e" => data <= x"0d";
            when "10" & x"e7f" => data <= x"6e";
            when "10" & x"e80" => data <= x"25";
            when "10" & x"e81" => data <= x"0d";
            when "10" & x"e82" => data <= x"6e";
            when "10" & x"e83" => data <= x"24";
            when "10" & x"e84" => data <= x"0d";
            when "10" & x"e85" => data <= x"6e";
            when "10" & x"e86" => data <= x"23";
            when "10" & x"e87" => data <= x"0d";
            when "10" & x"e88" => data <= x"20";
            when "10" & x"e89" => data <= x"a7";
            when "10" & x"e8a" => data <= x"aa";
            when "10" & x"e8b" => data <= x"38";
            when "10" & x"e8c" => data <= x"ad";
            when "10" & x"e8d" => data <= x"23";
            when "10" & x"e8e" => data <= x"0d";
            when "10" & x"e8f" => data <= x"09";
            when "10" & x"e90" => data <= x"0f";
            when "10" & x"e91" => data <= x"6d";
            when "10" & x"e92" => data <= x"06";
            when "10" & x"e93" => data <= x"0d";
            when "10" & x"e94" => data <= x"8d";
            when "10" & x"e95" => data <= x"23";
            when "10" & x"e96" => data <= x"0d";
            when "10" & x"e97" => data <= x"ad";
            when "10" & x"e98" => data <= x"24";
            when "10" & x"e99" => data <= x"0d";
            when "10" & x"e9a" => data <= x"6d";
            when "10" & x"e9b" => data <= x"07";
            when "10" & x"e9c" => data <= x"0d";
            when "10" & x"e9d" => data <= x"8d";
            when "10" & x"e9e" => data <= x"24";
            when "10" & x"e9f" => data <= x"0d";
            when "10" & x"ea0" => data <= x"ad";
            when "10" & x"ea1" => data <= x"25";
            when "10" & x"ea2" => data <= x"0d";
            when "10" & x"ea3" => data <= x"6d";
            when "10" & x"ea4" => data <= x"08";
            when "10" & x"ea5" => data <= x"0d";
            when "10" & x"ea6" => data <= x"8d";
            when "10" & x"ea7" => data <= x"25";
            when "10" & x"ea8" => data <= x"0d";
            when "10" & x"ea9" => data <= x"60";
            when "10" & x"eaa" => data <= x"a5";
            when "10" & x"eab" => data <= x"be";
            when "10" & x"eac" => data <= x"85";
            when "10" & x"ead" => data <= x"a0";
            when "10" & x"eae" => data <= x"a5";
            when "10" & x"eaf" => data <= x"bf";
            when "10" & x"eb0" => data <= x"85";
            when "10" & x"eb1" => data <= x"a1";
            when "10" & x"eb2" => data <= x"a6";
            when "10" & x"eb3" => data <= x"cf";
            when "10" & x"eb4" => data <= x"20";
            when "10" & x"eb5" => data <= x"1d";
            when "10" & x"eb6" => data <= x"ae";
            when "10" & x"eb7" => data <= x"18";
            when "10" & x"eb8" => data <= x"a5";
            when "10" & x"eb9" => data <= x"c4";
            when "10" & x"eba" => data <= x"29";
            when "10" & x"ebb" => data <= x"03";
            when "10" & x"ebc" => data <= x"48";
            when "10" & x"ebd" => data <= x"6a";
            when "10" & x"ebe" => data <= x"48";
            when "10" & x"ebf" => data <= x"a5";
            when "10" & x"ec0" => data <= x"c5";
            when "10" & x"ec1" => data <= x"6a";
            when "10" & x"ec2" => data <= x"48";
            when "10" & x"ec3" => data <= x"90";
            when "10" & x"ec4" => data <= x"03";
            when "10" & x"ec5" => data <= x"6e";
            when "10" & x"ec6" => data <= x"28";
            when "10" & x"ec7" => data <= x"0d";
            when "10" & x"ec8" => data <= x"18";
            when "10" & x"ec9" => data <= x"68";
            when "10" & x"eca" => data <= x"6d";
            when "10" & x"ecb" => data <= x"23";
            when "10" & x"ecc" => data <= x"0d";
            when "10" & x"ecd" => data <= x"8d";
            when "10" & x"ece" => data <= x"23";
            when "10" & x"ecf" => data <= x"0d";
            when "10" & x"ed0" => data <= x"68";
            when "10" & x"ed1" => data <= x"6d";
            when "10" & x"ed2" => data <= x"24";
            when "10" & x"ed3" => data <= x"0d";
            when "10" & x"ed4" => data <= x"8d";
            when "10" & x"ed5" => data <= x"24";
            when "10" & x"ed6" => data <= x"0d";
            when "10" & x"ed7" => data <= x"a9";
            when "10" & x"ed8" => data <= x"00";
            when "10" & x"ed9" => data <= x"6d";
            when "10" & x"eda" => data <= x"25";
            when "10" & x"edb" => data <= x"0d";
            when "10" & x"edc" => data <= x"8d";
            when "10" & x"edd" => data <= x"25";
            when "10" & x"ede" => data <= x"0d";
            when "10" & x"edf" => data <= x"a9";
            when "10" & x"ee0" => data <= x"00";
            when "10" & x"ee1" => data <= x"6d";
            when "10" & x"ee2" => data <= x"26";
            when "10" & x"ee3" => data <= x"0d";
            when "10" & x"ee4" => data <= x"8d";
            when "10" & x"ee5" => data <= x"26";
            when "10" & x"ee6" => data <= x"0d";
            when "10" & x"ee7" => data <= x"a5";
            when "10" & x"ee8" => data <= x"c3";
            when "10" & x"ee9" => data <= x"8d";
            when "10" & x"eea" => data <= x"27";
            when "10" & x"eeb" => data <= x"0d";
            when "10" & x"eec" => data <= x"a5";
            when "10" & x"eed" => data <= x"c4";
            when "10" & x"eee" => data <= x"4a";
            when "10" & x"eef" => data <= x"4a";
            when "10" & x"ef0" => data <= x"4a";
            when "10" & x"ef1" => data <= x"4a";
            when "10" & x"ef2" => data <= x"29";
            when "10" & x"ef3" => data <= x"03";
            when "10" & x"ef4" => data <= x"d0";
            when "10" & x"ef5" => data <= x"21";
            when "10" & x"ef6" => data <= x"a5";
            when "10" & x"ef7" => data <= x"c2";
            when "10" & x"ef8" => data <= x"8d";
            when "10" & x"ef9" => data <= x"29";
            when "10" & x"efa" => data <= x"0d";
            when "10" & x"efb" => data <= x"f0";
            when "10" & x"efc" => data <= x"05";
            when "10" & x"efd" => data <= x"ee";
            when "10" & x"efe" => data <= x"27";
            when "10" & x"eff" => data <= x"0d";
            when "10" & x"f00" => data <= x"f0";
            when "10" & x"f01" => data <= x"15";
            when "10" & x"f02" => data <= x"18";
            when "10" & x"f03" => data <= x"a5";
            when "10" & x"f04" => data <= x"c5";
            when "10" & x"f05" => data <= x"6d";
            when "10" & x"f06" => data <= x"27";
            when "10" & x"f07" => data <= x"0d";
            when "10" & x"f08" => data <= x"aa";
            when "10" & x"f09" => data <= x"68";
            when "10" & x"f0a" => data <= x"69";
            when "10" & x"f0b" => data <= x"00";
            when "10" & x"f0c" => data <= x"c9";
            when "10" & x"f0d" => data <= x"03";
            when "10" & x"f0e" => data <= x"90";
            when "10" & x"f0f" => data <= x"06";
            when "10" & x"f10" => data <= x"d0";
            when "10" & x"f11" => data <= x"17";
            when "10" & x"f12" => data <= x"e0";
            when "10" & x"f13" => data <= x"21";
            when "10" & x"f14" => data <= x"b0";
            when "10" & x"f15" => data <= x"13";
            when "10" & x"f16" => data <= x"60";
            when "10" & x"f17" => data <= x"20";
            when "10" & x"f18" => data <= x"00";
            when "10" & x"f19" => data <= x"a0";
            when "10" & x"f1a" => data <= x"ff";
            when "10" & x"f1b" => data <= x"42";
            when "10" & x"f1c" => data <= x"6c";
            when "10" & x"f1d" => data <= x"6f";
            when "10" & x"f1e" => data <= x"63";
            when "10" & x"f1f" => data <= x"6b";
            when "10" & x"f20" => data <= x"20";
            when "10" & x"f21" => data <= x"74";
            when "10" & x"f22" => data <= x"6f";
            when "10" & x"f23" => data <= x"6f";
            when "10" & x"f24" => data <= x"20";
            when "10" & x"f25" => data <= x"62";
            when "10" & x"f26" => data <= x"69";
            when "10" & x"f27" => data <= x"67";
            when "10" & x"f28" => data <= x"00";
            when "10" & x"f29" => data <= x"20";
            when "10" & x"f2a" => data <= x"00";
            when "10" & x"f2b" => data <= x"a0";
            when "10" & x"f2c" => data <= x"ff";
            when "10" & x"f2d" => data <= x"44";
            when "10" & x"f2e" => data <= x"69";
            when "10" & x"f2f" => data <= x"73";
            when "10" & x"f30" => data <= x"6b";
            when "10" & x"f31" => data <= x"20";
            when "10" & x"f32" => data <= x"6f";
            when "10" & x"f33" => data <= x"76";
            when "10" & x"f34" => data <= x"65";
            when "10" & x"f35" => data <= x"72";
            when "10" & x"f36" => data <= x"66";
            when "10" & x"f37" => data <= x"6c";
            when "10" & x"f38" => data <= x"6f";
            when "10" & x"f39" => data <= x"77";
            when "10" & x"f3a" => data <= x"00";
            when "10" & x"f3b" => data <= x"20";
            when "10" & x"f3c" => data <= x"4d";
            when "10" & x"f3d" => data <= x"83";
            when "10" & x"f3e" => data <= x"20";
            when "10" & x"f3f" => data <= x"58";
            when "10" & x"f40" => data <= x"83";
            when "10" & x"f41" => data <= x"20";
            when "10" & x"f42" => data <= x"1f";
            when "10" & x"f43" => data <= x"a6";
            when "10" & x"f44" => data <= x"a6";
            when "10" & x"f45" => data <= x"cf";
            when "10" & x"f46" => data <= x"8e";
            when "10" & x"f47" => data <= x"20";
            when "10" & x"f48" => data <= x"0d";
            when "10" & x"f49" => data <= x"20";
            when "10" & x"f4a" => data <= x"1d";
            when "10" & x"f4b" => data <= x"ae";
            when "10" & x"f4c" => data <= x"20";
            when "10" & x"f4d" => data <= x"99";
            when "10" & x"f4e" => data <= x"a7";
            when "10" & x"f4f" => data <= x"a5";
            when "10" & x"f50" => data <= x"cf";
            when "10" & x"f51" => data <= x"8d";
            when "10" & x"f52" => data <= x"82";
            when "10" & x"f53" => data <= x"10";
            when "10" & x"f54" => data <= x"60";
            when "10" & x"f55" => data <= x"20";
            when "10" & x"f56" => data <= x"1f";
            when "10" & x"f57" => data <= x"a6";
            when "10" & x"f58" => data <= x"a6";
            when "10" & x"f59" => data <= x"cf";
            when "10" & x"f5a" => data <= x"20";
            when "10" & x"f5b" => data <= x"cc";
            when "10" & x"f5c" => data <= x"ad";
            when "10" & x"f5d" => data <= x"20";
            when "10" & x"f5e" => data <= x"1d";
            when "10" & x"f5f" => data <= x"ae";
            when "10" & x"f60" => data <= x"4c";
            when "10" & x"f61" => data <= x"b2";
            when "10" & x"f62" => data <= x"a7";
            when "10" & x"f63" => data <= x"08";
            when "10" & x"f64" => data <= x"48";
            when "10" & x"f65" => data <= x"a0";
            when "10" & x"f66" => data <= x"ff";
            when "10" & x"f67" => data <= x"8c";
            when "10" & x"f68" => data <= x"82";
            when "10" & x"f69" => data <= x"10";
            when "10" & x"f6a" => data <= x"c8";
            when "10" & x"f6b" => data <= x"98";
            when "10" & x"f6c" => data <= x"99";
            when "10" & x"f6d" => data <= x"00";
            when "10" & x"f6e" => data <= x"0e";
            when "10" & x"f6f" => data <= x"99";
            when "10" & x"f70" => data <= x"00";
            when "10" & x"f71" => data <= x"0f";
            when "10" & x"f72" => data <= x"c8";
            when "10" & x"f73" => data <= x"d0";
            when "10" & x"f74" => data <= x"f7";
            when "10" & x"f75" => data <= x"a9";
            when "10" & x"f76" => data <= x"03";
            when "10" & x"f77" => data <= x"8d";
            when "10" & x"f78" => data <= x"06";
            when "10" & x"f79" => data <= x"0f";
            when "10" & x"f7a" => data <= x"a9";
            when "10" & x"f7b" => data <= x"20";
            when "10" & x"f7c" => data <= x"8d";
            when "10" & x"f7d" => data <= x"07";
            when "10" & x"f7e" => data <= x"0f";
            when "10" & x"f7f" => data <= x"20";
            when "10" & x"f80" => data <= x"1f";
            when "10" & x"f81" => data <= x"a6";
            when "10" & x"f82" => data <= x"68";
            when "10" & x"f83" => data <= x"28";
            when "10" & x"f84" => data <= x"20";
            when "10" & x"f85" => data <= x"26";
            when "10" & x"f86" => data <= x"ae";
            when "10" & x"f87" => data <= x"4c";
            when "10" & x"f88" => data <= x"b2";
            when "10" & x"f89" => data <= x"a7";
            when "10" & x"f8a" => data <= x"20";
            when "10" & x"f8b" => data <= x"1f";
            when "10" & x"f8c" => data <= x"a6";
            when "10" & x"f8d" => data <= x"20";
            when "10" & x"f8e" => data <= x"aa";
            when "10" & x"f8f" => data <= x"ae";
            when "10" & x"f90" => data <= x"20";
            when "10" & x"f91" => data <= x"cc";
            when "10" & x"f92" => data <= x"a7";
            when "10" & x"f93" => data <= x"20";
            when "10" & x"f94" => data <= x"cd";
            when "10" & x"f95" => data <= x"a0";
            when "10" & x"f96" => data <= x"a9";
            when "10" & x"f97" => data <= x"01";
            when "10" & x"f98" => data <= x"60";
            when "10" & x"f99" => data <= x"20";
            when "10" & x"f9a" => data <= x"1f";
            when "10" & x"f9b" => data <= x"a6";
            when "10" & x"f9c" => data <= x"20";
            when "10" & x"f9d" => data <= x"aa";
            when "10" & x"f9e" => data <= x"ae";
            when "10" & x"f9f" => data <= x"a6";
            when "10" & x"fa0" => data <= x"cf";
            when "10" & x"fa1" => data <= x"20";
            when "10" & x"fa2" => data <= x"cc";
            when "10" & x"fa3" => data <= x"ad";
            when "10" & x"fa4" => data <= x"20";
            when "10" & x"fa5" => data <= x"78";
            when "10" & x"fa6" => data <= x"a8";
            when "10" & x"fa7" => data <= x"20";
            when "10" & x"fa8" => data <= x"cd";
            when "10" & x"fa9" => data <= x"a0";
            when "10" & x"faa" => data <= x"a9";
            when "10" & x"fab" => data <= x"01";
            when "10" & x"fac" => data <= x"60";
            when "10" & x"fad" => data <= x"a8";
            when "10" & x"fae" => data <= x"c8";
            when "10" & x"faf" => data <= x"98";
            when "10" & x"fb0" => data <= x"d0";
            when "10" & x"fb1" => data <= x"01";
            when "10" & x"fb2" => data <= x"38";
            when "10" & x"fb3" => data <= x"2a";
            when "10" & x"fb4" => data <= x"2a";
            when "10" & x"fb5" => data <= x"2a";
            when "10" & x"fb6" => data <= x"2a";
            when "10" & x"fb7" => data <= x"2a";
            when "10" & x"fb8" => data <= x"48";
            when "10" & x"fb9" => data <= x"29";
            when "10" & x"fba" => data <= x"1f";
            when "10" & x"fbb" => data <= x"a8";
            when "10" & x"fbc" => data <= x"68";
            when "10" & x"fbd" => data <= x"09";
            when "10" & x"fbe" => data <= x"1f";
            when "10" & x"fbf" => data <= x"6a";
            when "10" & x"fc0" => data <= x"60";
            when "10" & x"fc1" => data <= x"20";
            when "10" & x"fc2" => data <= x"ad";
            when "10" & x"fc3" => data <= x"af";
            when "10" & x"fc4" => data <= x"48";
            when "10" & x"fc5" => data <= x"8a";
            when "10" & x"fc6" => data <= x"48";
            when "10" & x"fc7" => data <= x"98";
            when "10" & x"fc8" => data <= x"48";
            when "10" & x"fc9" => data <= x"20";
            when "10" & x"fca" => data <= x"97";
            when "10" & x"fcb" => data <= x"b0";
            when "10" & x"fcc" => data <= x"68";
            when "10" & x"fcd" => data <= x"6a";
            when "10" & x"fce" => data <= x"68";
            when "10" & x"fcf" => data <= x"aa";
            when "10" & x"fd0" => data <= x"68";
            when "10" & x"fd1" => data <= x"a8";
            when "10" & x"fd2" => data <= x"b0";
            when "10" & x"fd3" => data <= x"04";
            when "10" & x"fd4" => data <= x"b9";
            when "10" & x"fd5" => data <= x"00";
            when "10" & x"fd6" => data <= x"0e";
            when "10" & x"fd7" => data <= x"60";
            when "10" & x"fd8" => data <= x"b9";
            when "10" & x"fd9" => data <= x"00";
            when "10" & x"fda" => data <= x"0f";
            when "10" & x"fdb" => data <= x"60";
            when "10" & x"fdc" => data <= x"08";
            when "10" & x"fdd" => data <= x"48";
            when "10" & x"fde" => data <= x"8d";
            when "10" & x"fdf" => data <= x"5f";
            when "10" & x"fe0" => data <= x"0d";
            when "10" & x"fe1" => data <= x"a9";
            when "10" & x"fe2" => data <= x"00";
            when "10" & x"fe3" => data <= x"2a";
            when "10" & x"fe4" => data <= x"8d";
            when "10" & x"fe5" => data <= x"60";
            when "10" & x"fe6" => data <= x"0d";
            when "10" & x"fe7" => data <= x"8e";
            when "10" & x"fe8" => data <= x"61";
            when "10" & x"fe9" => data <= x"0d";
            when "10" & x"fea" => data <= x"a2";
            when "10" & x"feb" => data <= x"03";
            when "10" & x"fec" => data <= x"ec";
            when "10" & x"fed" => data <= x"61";
            when "10" & x"fee" => data <= x"0d";
            when "10" & x"fef" => data <= x"f0";
            when "10" & x"ff0" => data <= x"15";
            when "10" & x"ff1" => data <= x"bd";
            when "10" & x"ff2" => data <= x"0c";
            when "10" & x"ff3" => data <= x"0d";
            when "10" & x"ff4" => data <= x"cd";
            when "10" & x"ff5" => data <= x"5f";
            when "10" & x"ff6" => data <= x"0d";
            when "10" & x"ff7" => data <= x"d0";
            when "10" & x"ff8" => data <= x"0d";
            when "10" & x"ff9" => data <= x"bd";
            when "10" & x"ffa" => data <= x"10";
            when "10" & x"ffb" => data <= x"0d";
            when "10" & x"ffc" => data <= x"cd";
            when "10" & x"ffd" => data <= x"60";
            when "10" & x"ffe" => data <= x"0d";
            when "10" & x"fff" => data <= x"d0";
            when "11" & x"000" => data <= x"05";
            when "11" & x"001" => data <= x"a9";
            when "11" & x"002" => data <= x"ff";
            when "11" & x"003" => data <= x"9d";
            when "11" & x"004" => data <= x"10";
            when "11" & x"005" => data <= x"0d";
            when "11" & x"006" => data <= x"ca";
            when "11" & x"007" => data <= x"10";
            when "11" & x"008" => data <= x"e3";
            when "11" & x"009" => data <= x"ae";
            when "11" & x"00a" => data <= x"61";
            when "11" & x"00b" => data <= x"0d";
            when "11" & x"00c" => data <= x"68";
            when "11" & x"00d" => data <= x"28";
            when "11" & x"00e" => data <= x"60";
            when "11" & x"00f" => data <= x"08";
            when "11" & x"010" => data <= x"48";
            when "11" & x"011" => data <= x"9d";
            when "11" & x"012" => data <= x"0c";
            when "11" & x"013" => data <= x"0d";
            when "11" & x"014" => data <= x"49";
            when "11" & x"015" => data <= x"ff";
            when "11" & x"016" => data <= x"9d";
            when "11" & x"017" => data <= x"14";
            when "11" & x"018" => data <= x"0d";
            when "11" & x"019" => data <= x"a9";
            when "11" & x"01a" => data <= x"00";
            when "11" & x"01b" => data <= x"2a";
            when "11" & x"01c" => data <= x"9d";
            when "11" & x"01d" => data <= x"10";
            when "11" & x"01e" => data <= x"0d";
            when "11" & x"01f" => data <= x"49";
            when "11" & x"020" => data <= x"ff";
            when "11" & x"021" => data <= x"9d";
            when "11" & x"022" => data <= x"18";
            when "11" & x"023" => data <= x"0d";
            when "11" & x"024" => data <= x"68";
            when "11" & x"025" => data <= x"28";
            when "11" & x"026" => data <= x"20";
            when "11" & x"027" => data <= x"dc";
            when "11" & x"028" => data <= x"af";
            when "11" & x"029" => data <= x"20";
            when "11" & x"02a" => data <= x"c1";
            when "11" & x"02b" => data <= x"af";
            when "11" & x"02c" => data <= x"30";
            when "11" & x"02d" => data <= x"08";
            when "11" & x"02e" => data <= x"f0";
            when "11" & x"02f" => data <= x"03";
            when "11" & x"030" => data <= x"4c";
            when "11" & x"031" => data <= x"11";
            when "11" & x"032" => data <= x"ae";
            when "11" & x"033" => data <= x"4c";
            when "11" & x"034" => data <= x"17";
            when "11" & x"035" => data <= x"ae";
            when "11" & x"036" => data <= x"a8";
            when "11" & x"037" => data <= x"a9";
            when "11" & x"038" => data <= x"ff";
            when "11" & x"039" => data <= x"9d";
            when "11" & x"03a" => data <= x"10";
            when "11" & x"03b" => data <= x"0d";
            when "11" & x"03c" => data <= x"c8";
            when "11" & x"03d" => data <= x"d0";
            when "11" & x"03e" => data <= x"1a";
            when "11" & x"03f" => data <= x"20";
            when "11" & x"040" => data <= x"00";
            when "11" & x"041" => data <= x"a0";
            when "11" & x"042" => data <= x"c7";
            when "11" & x"043" => data <= x"44";
            when "11" & x"044" => data <= x"69";
            when "11" & x"045" => data <= x"73";
            when "11" & x"046" => data <= x"6b";
            when "11" & x"047" => data <= x"20";
            when "11" & x"048" => data <= x"6e";
            when "11" & x"049" => data <= x"75";
            when "11" & x"04a" => data <= x"6d";
            when "11" & x"04b" => data <= x"62";
            when "11" & x"04c" => data <= x"65";
            when "11" & x"04d" => data <= x"72";
            when "11" & x"04e" => data <= x"20";
            when "11" & x"04f" => data <= x"6e";
            when "11" & x"050" => data <= x"6f";
            when "11" & x"051" => data <= x"74";
            when "11" & x"052" => data <= x"20";
            when "11" & x"053" => data <= x"76";
            when "11" & x"054" => data <= x"61";
            when "11" & x"055" => data <= x"6c";
            when "11" & x"056" => data <= x"69";
            when "11" & x"057" => data <= x"64";
            when "11" & x"058" => data <= x"00";
            when "11" & x"059" => data <= x"20";
            when "11" & x"05a" => data <= x"00";
            when "11" & x"05b" => data <= x"a0";
            when "11" & x"05c" => data <= x"c7";
            when "11" & x"05d" => data <= x"44";
            when "11" & x"05e" => data <= x"69";
            when "11" & x"05f" => data <= x"73";
            when "11" & x"060" => data <= x"6b";
            when "11" & x"061" => data <= x"20";
            when "11" & x"062" => data <= x"6e";
            when "11" & x"063" => data <= x"6f";
            when "11" & x"064" => data <= x"74";
            when "11" & x"065" => data <= x"20";
            when "11" & x"066" => data <= x"66";
            when "11" & x"067" => data <= x"6f";
            when "11" & x"068" => data <= x"72";
            when "11" & x"069" => data <= x"6d";
            when "11" & x"06a" => data <= x"61";
            when "11" & x"06b" => data <= x"74";
            when "11" & x"06c" => data <= x"74";
            when "11" & x"06d" => data <= x"65";
            when "11" & x"06e" => data <= x"64";
            when "11" & x"06f" => data <= x"00";
            when "11" & x"070" => data <= x"29";
            when "11" & x"071" => data <= x"7f";
            when "11" & x"072" => data <= x"48";
            when "11" & x"073" => data <= x"20";
            when "11" & x"074" => data <= x"a7";
            when "11" & x"075" => data <= x"aa";
            when "11" & x"076" => data <= x"18";
            when "11" & x"077" => data <= x"68";
            when "11" & x"078" => data <= x"6d";
            when "11" & x"079" => data <= x"06";
            when "11" & x"07a" => data <= x"0d";
            when "11" & x"07b" => data <= x"8d";
            when "11" & x"07c" => data <= x"23";
            when "11" & x"07d" => data <= x"0d";
            when "11" & x"07e" => data <= x"ad";
            when "11" & x"07f" => data <= x"07";
            when "11" & x"080" => data <= x"0d";
            when "11" & x"081" => data <= x"69";
            when "11" & x"082" => data <= x"00";
            when "11" & x"083" => data <= x"8d";
            when "11" & x"084" => data <= x"24";
            when "11" & x"085" => data <= x"0d";
            when "11" & x"086" => data <= x"ad";
            when "11" & x"087" => data <= x"08";
            when "11" & x"088" => data <= x"0d";
            when "11" & x"089" => data <= x"69";
            when "11" & x"08a" => data <= x"00";
            when "11" & x"08b" => data <= x"8d";
            when "11" & x"08c" => data <= x"25";
            when "11" & x"08d" => data <= x"0d";
            when "11" & x"08e" => data <= x"ad";
            when "11" & x"08f" => data <= x"09";
            when "11" & x"090" => data <= x"0d";
            when "11" & x"091" => data <= x"69";
            when "11" & x"092" => data <= x"00";
            when "11" & x"093" => data <= x"8d";
            when "11" & x"094" => data <= x"26";
            when "11" & x"095" => data <= x"0d";
            when "11" & x"096" => data <= x"60";
            when "11" & x"097" => data <= x"29";
            when "11" & x"098" => data <= x"fe";
            when "11" & x"099" => data <= x"4a";
            when "11" & x"09a" => data <= x"09";
            when "11" & x"09b" => data <= x"80";
            when "11" & x"09c" => data <= x"cd";
            when "11" & x"09d" => data <= x"82";
            when "11" & x"09e" => data <= x"10";
            when "11" & x"09f" => data <= x"f0";
            when "11" & x"0a0" => data <= x"f5";
            when "11" & x"0a1" => data <= x"8d";
            when "11" & x"0a2" => data <= x"82";
            when "11" & x"0a3" => data <= x"10";
            when "11" & x"0a4" => data <= x"48";
            when "11" & x"0a5" => data <= x"20";
            when "11" & x"0a6" => data <= x"1f";
            when "11" & x"0a7" => data <= x"a6";
            when "11" & x"0a8" => data <= x"68";
            when "11" & x"0a9" => data <= x"20";
            when "11" & x"0aa" => data <= x"70";
            when "11" & x"0ab" => data <= x"b0";
            when "11" & x"0ac" => data <= x"4c";
            when "11" & x"0ad" => data <= x"99";
            when "11" & x"0ae" => data <= x"a7";
            when "11" & x"0af" => data <= x"8d";
            when "11" & x"0b0" => data <= x"82";
            when "11" & x"0b1" => data <= x"10";
            when "11" & x"0b2" => data <= x"20";
            when "11" & x"0b3" => data <= x"70";
            when "11" & x"0b4" => data <= x"b0";
            when "11" & x"0b5" => data <= x"4c";
            when "11" & x"0b6" => data <= x"99";
            when "11" & x"0b7" => data <= x"a7";
            when "11" & x"0b8" => data <= x"20";
            when "11" & x"0b9" => data <= x"1f";
            when "11" & x"0ba" => data <= x"a6";
            when "11" & x"0bb" => data <= x"ad";
            when "11" & x"0bc" => data <= x"82";
            when "11" & x"0bd" => data <= x"10";
            when "11" & x"0be" => data <= x"20";
            when "11" & x"0bf" => data <= x"70";
            when "11" & x"0c0" => data <= x"b0";
            when "11" & x"0c1" => data <= x"4c";
            when "11" & x"0c2" => data <= x"b2";
            when "11" & x"0c3" => data <= x"a7";
            when "11" & x"0c4" => data <= x"ad";
            when "11" & x"0c5" => data <= x"82";
            when "11" & x"0c6" => data <= x"10";
            when "11" & x"0c7" => data <= x"20";
            when "11" & x"0c8" => data <= x"70";
            when "11" & x"0c9" => data <= x"b0";
            when "11" & x"0ca" => data <= x"4c";
            when "11" & x"0cb" => data <= x"b2";
            when "11" & x"0cc" => data <= x"a7";
            when "11" & x"0cd" => data <= x"20";
            when "11" & x"0ce" => data <= x"b8";
            when "11" & x"0cf" => data <= x"b0";
            when "11" & x"0d0" => data <= x"a2";
            when "11" & x"0d1" => data <= x"03";
            when "11" & x"0d2" => data <= x"20";
            when "11" & x"0d3" => data <= x"d9";
            when "11" & x"0d4" => data <= x"b0";
            when "11" & x"0d5" => data <= x"ca";
            when "11" & x"0d6" => data <= x"10";
            when "11" & x"0d7" => data <= x"fa";
            when "11" & x"0d8" => data <= x"60";
            when "11" & x"0d9" => data <= x"bd";
            when "11" & x"0da" => data <= x"10";
            when "11" & x"0db" => data <= x"0d";
            when "11" & x"0dc" => data <= x"30";
            when "11" & x"0dd" => data <= x"2b";
            when "11" & x"0de" => data <= x"49";
            when "11" & x"0df" => data <= x"ff";
            when "11" & x"0e0" => data <= x"dd";
            when "11" & x"0e1" => data <= x"18";
            when "11" & x"0e2" => data <= x"0d";
            when "11" & x"0e3" => data <= x"d0";
            when "11" & x"0e4" => data <= x"18";
            when "11" & x"0e5" => data <= x"bd";
            when "11" & x"0e6" => data <= x"0c";
            when "11" & x"0e7" => data <= x"0d";
            when "11" & x"0e8" => data <= x"49";
            when "11" & x"0e9" => data <= x"ff";
            when "11" & x"0ea" => data <= x"dd";
            when "11" & x"0eb" => data <= x"14";
            when "11" & x"0ec" => data <= x"0d";
            when "11" & x"0ed" => data <= x"d0";
            when "11" & x"0ee" => data <= x"0e";
            when "11" & x"0ef" => data <= x"bd";
            when "11" & x"0f0" => data <= x"10";
            when "11" & x"0f1" => data <= x"0d";
            when "11" & x"0f2" => data <= x"6a";
            when "11" & x"0f3" => data <= x"bd";
            when "11" & x"0f4" => data <= x"0c";
            when "11" & x"0f5" => data <= x"0d";
            when "11" & x"0f6" => data <= x"20";
            when "11" & x"0f7" => data <= x"c1";
            when "11" & x"0f8" => data <= x"af";
            when "11" & x"0f9" => data <= x"f0";
            when "11" & x"0fa" => data <= x"0b";
            when "11" & x"0fb" => data <= x"10";
            when "11" & x"0fc" => data <= x"07";
            when "11" & x"0fd" => data <= x"a9";
            when "11" & x"0fe" => data <= x"ff";
            when "11" & x"0ff" => data <= x"9d";
            when "11" & x"100" => data <= x"10";
            when "11" & x"101" => data <= x"0d";
            when "11" & x"102" => data <= x"d0";
            when "11" & x"103" => data <= x"02";
            when "11" & x"104" => data <= x"a9";
            when "11" & x"105" => data <= x"54";
            when "11" & x"106" => data <= x"9d";
            when "11" & x"107" => data <= x"1c";
            when "11" & x"108" => data <= x"0d";
            when "11" & x"109" => data <= x"60";
            when "11" & x"10a" => data <= x"a2";
            when "11" & x"10b" => data <= x"00";
            when "11" & x"10c" => data <= x"bd";
            when "11" & x"10d" => data <= x"20";
            when "11" & x"10e" => data <= x"b3";
            when "11" & x"10f" => data <= x"9d";
            when "11" & x"110" => data <= x"70";
            when "11" & x"111" => data <= x"0d";
            when "11" & x"112" => data <= x"e8";
            when "11" & x"113" => data <= x"e0";
            when "11" & x"114" => data <= x"0b";
            when "11" & x"115" => data <= x"d0";
            when "11" & x"116" => data <= x"f5";
            when "11" & x"117" => data <= x"60";
            when "11" & x"118" => data <= x"a2";
            when "11" & x"119" => data <= x"6f";
            when "11" & x"11a" => data <= x"a9";
            when "11" & x"11b" => data <= x"00";
            when "11" & x"11c" => data <= x"9d";
            when "11" & x"11d" => data <= x"00";
            when "11" & x"11e" => data <= x"0d";
            when "11" & x"11f" => data <= x"ca";
            when "11" & x"120" => data <= x"d0";
            when "11" & x"121" => data <= x"fa";
            when "11" & x"122" => data <= x"a9";
            when "11" & x"123" => data <= x"40";
            when "11" & x"124" => data <= x"9d";
            when "11" & x"125" => data <= x"00";
            when "11" & x"126" => data <= x"0d";
            when "11" & x"127" => data <= x"60";
            when "11" & x"128" => data <= x"20";
            when "11" & x"129" => data <= x"0a";
            when "11" & x"12a" => data <= x"b1";
            when "11" & x"12b" => data <= x"20";
            when "11" & x"12c" => data <= x"18";
            when "11" & x"12d" => data <= x"b1";
            when "11" & x"12e" => data <= x"a9";
            when "11" & x"12f" => data <= x"ff";
            when "11" & x"130" => data <= x"8d";
            when "11" & x"131" => data <= x"52";
            when "11" & x"132" => data <= x"0d";
            when "11" & x"133" => data <= x"48";
            when "11" & x"134" => data <= x"4c";
            when "11" & x"135" => data <= x"3b";
            when "11" & x"136" => data <= x"93";
            when "11" & x"137" => data <= x"20";
            when "11" & x"138" => data <= x"0a";
            when "11" & x"139" => data <= x"b1";
            when "11" & x"13a" => data <= x"20";
            when "11" & x"13b" => data <= x"18";
            when "11" & x"13c" => data <= x"b1";
            when "11" & x"13d" => data <= x"a9";
            when "11" & x"13e" => data <= x"80";
            when "11" & x"13f" => data <= x"20";
            when "11" & x"140" => data <= x"a1";
            when "11" & x"141" => data <= x"b0";
            when "11" & x"142" => data <= x"a2";
            when "11" & x"143" => data <= x"00";
            when "11" & x"144" => data <= x"ad";
            when "11" & x"145" => data <= x"52";
            when "11" & x"146" => data <= x"0d";
            when "11" & x"147" => data <= x"c9";
            when "11" & x"148" => data <= x"42";
            when "11" & x"149" => data <= x"f0";
            when "11" & x"14a" => data <= x"16";
            when "11" & x"14b" => data <= x"bd";
            when "11" & x"14c" => data <= x"10";
            when "11" & x"14d" => data <= x"0d";
            when "11" & x"14e" => data <= x"30";
            when "11" & x"14f" => data <= x"43";
            when "11" & x"150" => data <= x"49";
            when "11" & x"151" => data <= x"ff";
            when "11" & x"152" => data <= x"dd";
            when "11" & x"153" => data <= x"18";
            when "11" & x"154" => data <= x"0d";
            when "11" & x"155" => data <= x"d0";
            when "11" & x"156" => data <= x"0a";
            when "11" & x"157" => data <= x"bd";
            when "11" & x"158" => data <= x"0c";
            when "11" & x"159" => data <= x"0d";
            when "11" & x"15a" => data <= x"49";
            when "11" & x"15b" => data <= x"ff";
            when "11" & x"15c" => data <= x"dd";
            when "11" & x"15d" => data <= x"14";
            when "11" & x"15e" => data <= x"0d";
            when "11" & x"15f" => data <= x"f0";
            when "11" & x"160" => data <= x"16";
            when "11" & x"161" => data <= x"bd";
            when "11" & x"162" => data <= x"00";
            when "11" & x"163" => data <= x"0e";
            when "11" & x"164" => data <= x"9d";
            when "11" & x"165" => data <= x"0c";
            when "11" & x"166" => data <= x"0d";
            when "11" & x"167" => data <= x"49";
            when "11" & x"168" => data <= x"ff";
            when "11" & x"169" => data <= x"9d";
            when "11" & x"16a" => data <= x"14";
            when "11" & x"16b" => data <= x"0d";
            when "11" & x"16c" => data <= x"bd";
            when "11" & x"16d" => data <= x"04";
            when "11" & x"16e" => data <= x"0e";
            when "11" & x"16f" => data <= x"9d";
            when "11" & x"170" => data <= x"10";
            when "11" & x"171" => data <= x"0d";
            when "11" & x"172" => data <= x"49";
            when "11" & x"173" => data <= x"ff";
            when "11" & x"174" => data <= x"9d";
            when "11" & x"175" => data <= x"18";
            when "11" & x"176" => data <= x"0d";
            when "11" & x"177" => data <= x"8a";
            when "11" & x"178" => data <= x"f0";
            when "11" & x"179" => data <= x"1e";
            when "11" & x"17a" => data <= x"a8";
            when "11" & x"17b" => data <= x"88";
            when "11" & x"17c" => data <= x"bd";
            when "11" & x"17d" => data <= x"10";
            when "11" & x"17e" => data <= x"0d";
            when "11" & x"17f" => data <= x"30";
            when "11" & x"180" => data <= x"17";
            when "11" & x"181" => data <= x"d9";
            when "11" & x"182" => data <= x"10";
            when "11" & x"183" => data <= x"0d";
            when "11" & x"184" => data <= x"d0";
            when "11" & x"185" => data <= x"08";
            when "11" & x"186" => data <= x"bd";
            when "11" & x"187" => data <= x"0c";
            when "11" & x"188" => data <= x"0d";
            when "11" & x"189" => data <= x"d9";
            when "11" & x"18a" => data <= x"0c";
            when "11" & x"18b" => data <= x"0d";
            when "11" & x"18c" => data <= x"f0";
            when "11" & x"18d" => data <= x"05";
            when "11" & x"18e" => data <= x"88";
            when "11" & x"18f" => data <= x"10";
            when "11" & x"190" => data <= x"eb";
            when "11" & x"191" => data <= x"30";
            when "11" & x"192" => data <= x"05";
            when "11" & x"193" => data <= x"a9";
            when "11" & x"194" => data <= x"ff";
            when "11" & x"195" => data <= x"9d";
            when "11" & x"196" => data <= x"10";
            when "11" & x"197" => data <= x"0d";
            when "11" & x"198" => data <= x"e8";
            when "11" & x"199" => data <= x"e0";
            when "11" & x"19a" => data <= x"04";
            when "11" & x"19b" => data <= x"d0";
            when "11" & x"19c" => data <= x"a7";
            when "11" & x"19d" => data <= x"4c";
            when "11" & x"19e" => data <= x"d0";
            when "11" & x"19f" => data <= x"b0";
            when "11" & x"1a0" => data <= x"08";
            when "11" & x"1a1" => data <= x"48";
            when "11" & x"1a2" => data <= x"8d";
            when "11" & x"1a3" => data <= x"53";
            when "11" & x"1a4" => data <= x"0d";
            when "11" & x"1a5" => data <= x"a9";
            when "11" & x"1a6" => data <= x"00";
            when "11" & x"1a7" => data <= x"2a";
            when "11" & x"1a8" => data <= x"8d";
            when "11" & x"1a9" => data <= x"54";
            when "11" & x"1aa" => data <= x"0d";
            when "11" & x"1ab" => data <= x"68";
            when "11" & x"1ac" => data <= x"28";
            when "11" & x"1ad" => data <= x"08";
            when "11" & x"1ae" => data <= x"48";
            when "11" & x"1af" => data <= x"20";
            when "11" & x"1b0" => data <= x"6c";
            when "11" & x"1b1" => data <= x"ad";
            when "11" & x"1b2" => data <= x"8e";
            when "11" & x"1b3" => data <= x"55";
            when "11" & x"1b4" => data <= x"0d";
            when "11" & x"1b5" => data <= x"8d";
            when "11" & x"1b6" => data <= x"56";
            when "11" & x"1b7" => data <= x"0d";
            when "11" & x"1b8" => data <= x"68";
            when "11" & x"1b9" => data <= x"28";
            when "11" & x"1ba" => data <= x"20";
            when "11" & x"1bb" => data <= x"ad";
            when "11" & x"1bc" => data <= x"af";
            when "11" & x"1bd" => data <= x"29";
            when "11" & x"1be" => data <= x"f0";
            when "11" & x"1bf" => data <= x"85";
            when "11" & x"1c0" => data <= x"f2";
            when "11" & x"1c1" => data <= x"98";
            when "11" & x"1c2" => data <= x"29";
            when "11" & x"1c3" => data <= x"01";
            when "11" & x"1c4" => data <= x"09";
            when "11" & x"1c5" => data <= x"0e";
            when "11" & x"1c6" => data <= x"85";
            when "11" & x"1c7" => data <= x"f3";
            when "11" & x"1c8" => data <= x"98";
            when "11" & x"1c9" => data <= x"29";
            when "11" & x"1ca" => data <= x"fe";
            when "11" & x"1cb" => data <= x"4a";
            when "11" & x"1cc" => data <= x"09";
            when "11" & x"1cd" => data <= x"80";
            when "11" & x"1ce" => data <= x"8d";
            when "11" & x"1cf" => data <= x"52";
            when "11" & x"1d0" => data <= x"0d";
            when "11" & x"1d1" => data <= x"20";
            when "11" & x"1d2" => data <= x"9c";
            when "11" & x"1d3" => data <= x"b0";
            when "11" & x"1d4" => data <= x"4c";
            when "11" & x"1d5" => data <= x"35";
            when "11" & x"1d6" => data <= x"b2";
            when "11" & x"1d7" => data <= x"a9";
            when "11" & x"1d8" => data <= x"00";
            when "11" & x"1d9" => data <= x"8d";
            when "11" & x"1da" => data <= x"55";
            when "11" & x"1db" => data <= x"0d";
            when "11" & x"1dc" => data <= x"8d";
            when "11" & x"1dd" => data <= x"56";
            when "11" & x"1de" => data <= x"0d";
            when "11" & x"1df" => data <= x"8d";
            when "11" & x"1e0" => data <= x"53";
            when "11" & x"1e1" => data <= x"0d";
            when "11" & x"1e2" => data <= x"8d";
            when "11" & x"1e3" => data <= x"54";
            when "11" & x"1e4" => data <= x"0d";
            when "11" & x"1e5" => data <= x"a9";
            when "11" & x"1e6" => data <= x"10";
            when "11" & x"1e7" => data <= x"85";
            when "11" & x"1e8" => data <= x"f2";
            when "11" & x"1e9" => data <= x"a9";
            when "11" & x"1ea" => data <= x"0e";
            when "11" & x"1eb" => data <= x"85";
            when "11" & x"1ec" => data <= x"f3";
            when "11" & x"1ed" => data <= x"a9";
            when "11" & x"1ee" => data <= x"80";
            when "11" & x"1ef" => data <= x"8d";
            when "11" & x"1f0" => data <= x"52";
            when "11" & x"1f1" => data <= x"0d";
            when "11" & x"1f2" => data <= x"20";
            when "11" & x"1f3" => data <= x"9c";
            when "11" & x"1f4" => data <= x"b0";
            when "11" & x"1f5" => data <= x"4c";
            when "11" & x"1f6" => data <= x"35";
            when "11" & x"1f7" => data <= x"b2";
            when "11" & x"1f8" => data <= x"c9";
            when "11" & x"1f9" => data <= x"ff";
            when "11" & x"1fa" => data <= x"f0";
            when "11" & x"1fb" => data <= x"41";
            when "11" & x"1fc" => data <= x"18";
            when "11" & x"1fd" => data <= x"a5";
            when "11" & x"1fe" => data <= x"f2";
            when "11" & x"1ff" => data <= x"69";
            when "11" & x"200" => data <= x"10";
            when "11" & x"201" => data <= x"85";
            when "11" & x"202" => data <= x"f2";
            when "11" & x"203" => data <= x"d0";
            when "11" & x"204" => data <= x"18";
            when "11" & x"205" => data <= x"a5";
            when "11" & x"206" => data <= x"f3";
            when "11" & x"207" => data <= x"49";
            when "11" & x"208" => data <= x"01";
            when "11" & x"209" => data <= x"85";
            when "11" & x"20a" => data <= x"f3";
            when "11" & x"20b" => data <= x"6a";
            when "11" & x"20c" => data <= x"b0";
            when "11" & x"20d" => data <= x"0f";
            when "11" & x"20e" => data <= x"ad";
            when "11" & x"20f" => data <= x"52";
            when "11" & x"210" => data <= x"0d";
            when "11" & x"211" => data <= x"69";
            when "11" & x"212" => data <= x"01";
            when "11" & x"213" => data <= x"c9";
            when "11" & x"214" => data <= x"90";
            when "11" & x"215" => data <= x"f0";
            when "11" & x"216" => data <= x"26";
            when "11" & x"217" => data <= x"8d";
            when "11" & x"218" => data <= x"52";
            when "11" & x"219" => data <= x"0d";
            when "11" & x"21a" => data <= x"20";
            when "11" & x"21b" => data <= x"9c";
            when "11" & x"21c" => data <= x"b0";
            when "11" & x"21d" => data <= x"ee";
            when "11" & x"21e" => data <= x"53";
            when "11" & x"21f" => data <= x"0d";
            when "11" & x"220" => data <= x"d0";
            when "11" & x"221" => data <= x"03";
            when "11" & x"222" => data <= x"ee";
            when "11" & x"223" => data <= x"54";
            when "11" & x"224" => data <= x"0d";
            when "11" & x"225" => data <= x"f8";
            when "11" & x"226" => data <= x"18";
            when "11" & x"227" => data <= x"ad";
            when "11" & x"228" => data <= x"55";
            when "11" & x"229" => data <= x"0d";
            when "11" & x"22a" => data <= x"69";
            when "11" & x"22b" => data <= x"01";
            when "11" & x"22c" => data <= x"8d";
            when "11" & x"22d" => data <= x"55";
            when "11" & x"22e" => data <= x"0d";
            when "11" & x"22f" => data <= x"90";
            when "11" & x"230" => data <= x"03";
            when "11" & x"231" => data <= x"ee";
            when "11" & x"232" => data <= x"56";
            when "11" & x"233" => data <= x"0d";
            when "11" & x"234" => data <= x"d8";
            when "11" & x"235" => data <= x"a0";
            when "11" & x"236" => data <= x"0f";
            when "11" & x"237" => data <= x"b1";
            when "11" & x"238" => data <= x"f2";
            when "11" & x"239" => data <= x"30";
            when "11" & x"23a" => data <= x"bd";
            when "11" & x"23b" => data <= x"18";
            when "11" & x"23c" => data <= x"60";
            when "11" & x"23d" => data <= x"a9";
            when "11" & x"23e" => data <= x"ff";
            when "11" & x"23f" => data <= x"8d";
            when "11" & x"240" => data <= x"54";
            when "11" & x"241" => data <= x"0d";
            when "11" & x"242" => data <= x"38";
            when "11" & x"243" => data <= x"60";
            when "11" & x"244" => data <= x"20";
            when "11" & x"245" => data <= x"1f";
            when "11" & x"246" => data <= x"a6";
            when "11" & x"247" => data <= x"a9";
            when "11" & x"248" => data <= x"80";
            when "11" & x"249" => data <= x"8d";
            when "11" & x"24a" => data <= x"52";
            when "11" & x"24b" => data <= x"0d";
            when "11" & x"24c" => data <= x"20";
            when "11" & x"24d" => data <= x"af";
            when "11" & x"24e" => data <= x"b0";
            when "11" & x"24f" => data <= x"a9";
            when "11" & x"250" => data <= x"10";
            when "11" & x"251" => data <= x"85";
            when "11" & x"252" => data <= x"f2";
            when "11" & x"253" => data <= x"a9";
            when "11" & x"254" => data <= x"0e";
            when "11" & x"255" => data <= x"85";
            when "11" & x"256" => data <= x"f3";
            when "11" & x"257" => data <= x"20";
            when "11" & x"258" => data <= x"a7";
            when "11" & x"259" => data <= x"aa";
            when "11" & x"25a" => data <= x"18";
            when "11" & x"25b" => data <= x"ad";
            when "11" & x"25c" => data <= x"06";
            when "11" & x"25d" => data <= x"0d";
            when "11" & x"25e" => data <= x"69";
            when "11" & x"25f" => data <= x"10";
            when "11" & x"260" => data <= x"8d";
            when "11" & x"261" => data <= x"23";
            when "11" & x"262" => data <= x"0d";
            when "11" & x"263" => data <= x"ad";
            when "11" & x"264" => data <= x"07";
            when "11" & x"265" => data <= x"0d";
            when "11" & x"266" => data <= x"69";
            when "11" & x"267" => data <= x"00";
            when "11" & x"268" => data <= x"8d";
            when "11" & x"269" => data <= x"24";
            when "11" & x"26a" => data <= x"0d";
            when "11" & x"26b" => data <= x"ad";
            when "11" & x"26c" => data <= x"08";
            when "11" & x"26d" => data <= x"0d";
            when "11" & x"26e" => data <= x"69";
            when "11" & x"26f" => data <= x"00";
            when "11" & x"270" => data <= x"8d";
            when "11" & x"271" => data <= x"25";
            when "11" & x"272" => data <= x"0d";
            when "11" & x"273" => data <= x"ad";
            when "11" & x"274" => data <= x"09";
            when "11" & x"275" => data <= x"0d";
            when "11" & x"276" => data <= x"69";
            when "11" & x"277" => data <= x"00";
            when "11" & x"278" => data <= x"8d";
            when "11" & x"279" => data <= x"09";
            when "11" & x"27a" => data <= x"0d";
            when "11" & x"27b" => data <= x"20";
            when "11" & x"27c" => data <= x"1e";
            when "11" & x"27d" => data <= x"a9";
            when "11" & x"27e" => data <= x"a0";
            when "11" & x"27f" => data <= x"0f";
            when "11" & x"280" => data <= x"b1";
            when "11" & x"281" => data <= x"f2";
            when "11" & x"282" => data <= x"c9";
            when "11" & x"283" => data <= x"ff";
            when "11" & x"284" => data <= x"f0";
            when "11" & x"285" => data <= x"39";
            when "11" & x"286" => data <= x"20";
            when "11" & x"287" => data <= x"24";
            when "11" & x"288" => data <= x"a9";
            when "11" & x"289" => data <= x"a0";
            when "11" & x"28a" => data <= x"0b";
            when "11" & x"28b" => data <= x"b9";
            when "11" & x"28c" => data <= x"5f";
            when "11" & x"28d" => data <= x"0d";
            when "11" & x"28e" => data <= x"91";
            when "11" & x"28f" => data <= x"f2";
            when "11" & x"290" => data <= x"88";
            when "11" & x"291" => data <= x"10";
            when "11" & x"292" => data <= x"f8";
            when "11" & x"293" => data <= x"18";
            when "11" & x"294" => data <= x"a5";
            when "11" & x"295" => data <= x"f2";
            when "11" & x"296" => data <= x"69";
            when "11" & x"297" => data <= x"10";
            when "11" & x"298" => data <= x"85";
            when "11" & x"299" => data <= x"f2";
            when "11" & x"29a" => data <= x"d0";
            when "11" & x"29b" => data <= x"e2";
            when "11" & x"29c" => data <= x"a5";
            when "11" & x"29d" => data <= x"f3";
            when "11" & x"29e" => data <= x"49";
            when "11" & x"29f" => data <= x"01";
            when "11" & x"2a0" => data <= x"85";
            when "11" & x"2a1" => data <= x"f3";
            when "11" & x"2a2" => data <= x"6a";
            when "11" & x"2a3" => data <= x"b0";
            when "11" & x"2a4" => data <= x"d9";
            when "11" & x"2a5" => data <= x"20";
            when "11" & x"2a6" => data <= x"c4";
            when "11" & x"2a7" => data <= x"b0";
            when "11" & x"2a8" => data <= x"18";
            when "11" & x"2a9" => data <= x"ad";
            when "11" & x"2aa" => data <= x"52";
            when "11" & x"2ab" => data <= x"0d";
            when "11" & x"2ac" => data <= x"69";
            when "11" & x"2ad" => data <= x"01";
            when "11" & x"2ae" => data <= x"c9";
            when "11" & x"2af" => data <= x"90";
            when "11" & x"2b0" => data <= x"f0";
            when "11" & x"2b1" => data <= x"18";
            when "11" & x"2b2" => data <= x"8d";
            when "11" & x"2b3" => data <= x"52";
            when "11" & x"2b4" => data <= x"0d";
            when "11" & x"2b5" => data <= x"24";
            when "11" & x"2b6" => data <= x"ff";
            when "11" & x"2b7" => data <= x"30";
            when "11" & x"2b8" => data <= x"12";
            when "11" & x"2b9" => data <= x"20";
            when "11" & x"2ba" => data <= x"af";
            when "11" & x"2bb" => data <= x"b0";
            when "11" & x"2bc" => data <= x"4c";
            when "11" & x"2bd" => data <= x"7e";
            when "11" & x"2be" => data <= x"b2";
            when "11" & x"2bf" => data <= x"a5";
            when "11" & x"2c0" => data <= x"f2";
            when "11" & x"2c1" => data <= x"d0";
            when "11" & x"2c2" => data <= x"04";
            when "11" & x"2c3" => data <= x"66";
            when "11" & x"2c4" => data <= x"f3";
            when "11" & x"2c5" => data <= x"90";
            when "11" & x"2c6" => data <= x"03";
            when "11" & x"2c7" => data <= x"20";
            when "11" & x"2c8" => data <= x"c4";
            when "11" & x"2c9" => data <= x"b0";
            when "11" & x"2ca" => data <= x"60";
            when "11" & x"2cb" => data <= x"4c";
            when "11" & x"2cc" => data <= x"82";
            when "11" & x"2cd" => data <= x"a0";
            when "11" & x"2ce" => data <= x"a2";
            when "11" & x"2cf" => data <= x"0b";
            when "11" & x"2d0" => data <= x"a9";
            when "11" & x"2d1" => data <= x"00";
            when "11" & x"2d2" => data <= x"20";
            when "11" & x"2d3" => data <= x"c6";
            when "11" & x"2d4" => data <= x"88";
            when "11" & x"2d5" => data <= x"9d";
            when "11" & x"2d6" => data <= x"5f";
            when "11" & x"2d7" => data <= x"0d";
            when "11" & x"2d8" => data <= x"ca";
            when "11" & x"2d9" => data <= x"10";
            when "11" & x"2da" => data <= x"f7";
            when "11" & x"2db" => data <= x"e8";
            when "11" & x"2dc" => data <= x"20";
            when "11" & x"2dd" => data <= x"c5";
            when "11" & x"2de" => data <= x"ff";
            when "11" & x"2df" => data <= x"b0";
            when "11" & x"2e0" => data <= x"0a";
            when "11" & x"2e1" => data <= x"20";
            when "11" & x"2e2" => data <= x"c6";
            when "11" & x"2e3" => data <= x"88";
            when "11" & x"2e4" => data <= x"9d";
            when "11" & x"2e5" => data <= x"5f";
            when "11" & x"2e6" => data <= x"0d";
            when "11" & x"2e7" => data <= x"e0";
            when "11" & x"2e8" => data <= x"0b";
            when "11" & x"2e9" => data <= x"90";
            when "11" & x"2ea" => data <= x"f0";
            when "11" & x"2eb" => data <= x"20";
            when "11" & x"2ec" => data <= x"b4";
            when "11" & x"2ed" => data <= x"8a";
            when "11" & x"2ee" => data <= x"ae";
            when "11" & x"2ef" => data <= x"82";
            when "11" & x"2f0" => data <= x"10";
            when "11" & x"2f1" => data <= x"bd";
            when "11" & x"2f2" => data <= x"10";
            when "11" & x"2f3" => data <= x"0d";
            when "11" & x"2f4" => data <= x"6a";
            when "11" & x"2f5" => data <= x"bd";
            when "11" & x"2f6" => data <= x"0c";
            when "11" & x"2f7" => data <= x"0d";
            when "11" & x"2f8" => data <= x"20";
            when "11" & x"2f9" => data <= x"ad";
            when "11" & x"2fa" => data <= x"af";
            when "11" & x"2fb" => data <= x"29";
            when "11" & x"2fc" => data <= x"f0";
            when "11" & x"2fd" => data <= x"48";
            when "11" & x"2fe" => data <= x"98";
            when "11" & x"2ff" => data <= x"48";
            when "11" & x"300" => data <= x"29";
            when "11" & x"301" => data <= x"fe";
            when "11" & x"302" => data <= x"4a";
            when "11" & x"303" => data <= x"09";
            when "11" & x"304" => data <= x"80";
            when "11" & x"305" => data <= x"20";
            when "11" & x"306" => data <= x"a1";
            when "11" & x"307" => data <= x"b0";
            when "11" & x"308" => data <= x"68";
            when "11" & x"309" => data <= x"18";
            when "11" & x"30a" => data <= x"29";
            when "11" & x"30b" => data <= x"01";
            when "11" & x"30c" => data <= x"69";
            when "11" & x"30d" => data <= x"0e";
            when "11" & x"30e" => data <= x"85";
            when "11" & x"30f" => data <= x"f3";
            when "11" & x"310" => data <= x"68";
            when "11" & x"311" => data <= x"85";
            when "11" & x"312" => data <= x"f2";
            when "11" & x"313" => data <= x"a0";
            when "11" & x"314" => data <= x"0b";
            when "11" & x"315" => data <= x"b9";
            when "11" & x"316" => data <= x"5f";
            when "11" & x"317" => data <= x"0d";
            when "11" & x"318" => data <= x"91";
            when "11" & x"319" => data <= x"f2";
            when "11" & x"31a" => data <= x"88";
            when "11" & x"31b" => data <= x"10";
            when "11" & x"31c" => data <= x"f8";
            when "11" & x"31d" => data <= x"4c";
            when "11" & x"31e" => data <= x"b8";
            when "11" & x"31f" => data <= x"b0";
            when "11" & x"320" => data <= x"42";
            when "11" & x"321" => data <= x"45";
            when "11" & x"322" => data <= x"45";
            when "11" & x"323" => data <= x"42";
            when "11" & x"324" => data <= x"20";
            when "11" & x"325" => data <= x"20";
            when "11" & x"326" => data <= x"20";
            when "11" & x"327" => data <= x"20";
            when "11" & x"328" => data <= x"4d";
            when "11" & x"329" => data <= x"4d";
            when "11" & x"32a" => data <= x"42";
            when "11" & x"32b" => data <= x"44";
            when "11" & x"32c" => data <= x"49";
            when "11" & x"32d" => data <= x"4e";
            when "11" & x"32e" => data <= x"b8";
            when "11" & x"32f" => data <= x"05";
            when "11" & x"330" => data <= x"12";
            when "11" & x"331" => data <= x"44";
            when "11" & x"332" => data <= x"42";
            when "11" & x"333" => data <= x"4f";
            when "11" & x"334" => data <= x"4f";
            when "11" & x"335" => data <= x"54";
            when "11" & x"336" => data <= x"b7";
            when "11" & x"337" => data <= x"fa";
            when "11" & x"338" => data <= x"02";
            when "11" & x"339" => data <= x"44";
            when "11" & x"33a" => data <= x"43";
            when "11" & x"33b" => data <= x"41";
            when "11" & x"33c" => data <= x"54";
            when "11" & x"33d" => data <= x"b8";
            when "11" & x"33e" => data <= x"0b";
            when "11" & x"33f" => data <= x"04";
            when "11" & x"340" => data <= x"44";
            when "11" & x"341" => data <= x"44";
            when "11" & x"342" => data <= x"49";
            when "11" & x"343" => data <= x"53";
            when "11" & x"344" => data <= x"4b";
            when "11" & x"345" => data <= x"53";
            when "11" & x"346" => data <= x"b9";
            when "11" & x"347" => data <= x"bb";
            when "11" & x"348" => data <= x"01";
            when "11" & x"349" => data <= x"44";
            when "11" & x"34a" => data <= x"4c";
            when "11" & x"34b" => data <= x"4f";
            when "11" & x"34c" => data <= x"43";
            when "11" & x"34d" => data <= x"4b";
            when "11" & x"34e" => data <= x"ba";
            when "11" & x"34f" => data <= x"01";
            when "11" & x"350" => data <= x"02";
            when "11" & x"351" => data <= x"44";
            when "11" & x"352" => data <= x"55";
            when "11" & x"353" => data <= x"4e";
            when "11" & x"354" => data <= x"4c";
            when "11" & x"355" => data <= x"4f";
            when "11" & x"356" => data <= x"43";
            when "11" & x"357" => data <= x"4b";
            when "11" & x"358" => data <= x"ba";
            when "11" & x"359" => data <= x"05";
            when "11" & x"35a" => data <= x"02";
            when "11" & x"35b" => data <= x"44";
            when "11" & x"35c" => data <= x"46";
            when "11" & x"35d" => data <= x"52";
            when "11" & x"35e" => data <= x"45";
            when "11" & x"35f" => data <= x"45";
            when "11" & x"360" => data <= x"b8";
            when "11" & x"361" => data <= x"f5";
            when "11" & x"362" => data <= x"00";
            when "11" & x"363" => data <= x"44";
            when "11" & x"364" => data <= x"4b";
            when "11" & x"365" => data <= x"49";
            when "11" & x"366" => data <= x"4c";
            when "11" & x"367" => data <= x"4c";
            when "11" & x"368" => data <= x"ba";
            when "11" & x"369" => data <= x"28";
            when "11" & x"36a" => data <= x"03";
            when "11" & x"36b" => data <= x"44";
            when "11" & x"36c" => data <= x"52";
            when "11" & x"36d" => data <= x"45";
            when "11" & x"36e" => data <= x"53";
            when "11" & x"36f" => data <= x"54";
            when "11" & x"370" => data <= x"4f";
            when "11" & x"371" => data <= x"52";
            when "11" & x"372" => data <= x"45";
            when "11" & x"373" => data <= x"ba";
            when "11" & x"374" => data <= x"6b";
            when "11" & x"375" => data <= x"03";
            when "11" & x"376" => data <= x"44";
            when "11" & x"377" => data <= x"4e";
            when "11" & x"378" => data <= x"45";
            when "11" & x"379" => data <= x"57";
            when "11" & x"37a" => data <= x"ba";
            when "11" & x"37b" => data <= x"c0";
            when "11" & x"37c" => data <= x"01";
            when "11" & x"37d" => data <= x"44";
            when "11" & x"37e" => data <= x"46";
            when "11" & x"37f" => data <= x"4f";
            when "11" & x"380" => data <= x"52";
            when "11" & x"381" => data <= x"4d";
            when "11" & x"382" => data <= x"ba";
            when "11" & x"383" => data <= x"63";
            when "11" & x"384" => data <= x"03";
            when "11" & x"385" => data <= x"44";
            when "11" & x"386" => data <= x"4f";
            when "11" & x"387" => data <= x"4e";
            when "11" & x"388" => data <= x"42";
            when "11" & x"389" => data <= x"4f";
            when "11" & x"38a" => data <= x"4f";
            when "11" & x"38b" => data <= x"54";
            when "11" & x"38c" => data <= x"bb";
            when "11" & x"38d" => data <= x"8e";
            when "11" & x"38e" => data <= x"52";
            when "11" & x"38f" => data <= x"44";
            when "11" & x"390" => data <= x"52";
            when "11" & x"391" => data <= x"45";
            when "11" & x"392" => data <= x"43";
            when "11" & x"393" => data <= x"41";
            when "11" & x"394" => data <= x"54";
            when "11" & x"395" => data <= x"b2";
            when "11" & x"396" => data <= x"43";
            when "11" & x"397" => data <= x"00";
            when "11" & x"398" => data <= x"44";
            when "11" & x"399" => data <= x"52";
            when "11" & x"39a" => data <= x"4f";
            when "11" & x"39b" => data <= x"4d";
            when "11" & x"39c" => data <= x"bc";
            when "11" & x"39d" => data <= x"1a";
            when "11" & x"39e" => data <= x"86";
            when "11" & x"39f" => data <= x"42";
            when "11" & x"3a0" => data <= x"45";
            when "11" & x"3a1" => data <= x"45";
            when "11" & x"3a2" => data <= x"42";
            when "11" & x"3a3" => data <= x"bb";
            when "11" & x"3a4" => data <= x"a9";
            when "11" & x"3a5" => data <= x"03";
            when "11" & x"3a6" => data <= x"44";
            when "11" & x"3a7" => data <= x"47";
            when "11" & x"3a8" => data <= x"45";
            when "11" & x"3a9" => data <= x"54";
            when "11" & x"3aa" => data <= x"bc";
            when "11" & x"3ab" => data <= x"14";
            when "11" & x"3ac" => data <= x"00";
            when "11" & x"3ad" => data <= x"44";
            when "11" & x"3ae" => data <= x"50";
            when "11" & x"3af" => data <= x"55";
            when "11" & x"3b0" => data <= x"54";
            when "11" & x"3b1" => data <= x"bc";
            when "11" & x"3b2" => data <= x"17";
            when "11" & x"3b3" => data <= x"00";
            when "11" & x"3b4" => data <= x"44";
            when "11" & x"3b5" => data <= x"41";
            when "11" & x"3b6" => data <= x"42";
            when "11" & x"3b7" => data <= x"4f";
            when "11" & x"3b8" => data <= x"55";
            when "11" & x"3b9" => data <= x"54";
            when "11" & x"3ba" => data <= x"b4";
            when "11" & x"3bb" => data <= x"32";
            when "11" & x"3bc" => data <= x"00";
            when "11" & x"3bd" => data <= x"87";
            when "11" & x"3be" => data <= x"d6";
            when "11" & x"3bf" => data <= x"00";
            when "11" & x"3c0" => data <= x"44";
            when "11" & x"3c1" => data <= x"55";
            when "11" & x"3c2" => data <= x"54";
            when "11" & x"3c3" => data <= x"49";
            when "11" & x"3c4" => data <= x"4c";
            when "11" & x"3c5" => data <= x"53";
            when "11" & x"3c6" => data <= x"b4";
            when "11" & x"3c7" => data <= x"03";
            when "11" & x"3c8" => data <= x"00";
            when "11" & x"3c9" => data <= x"b3";
            when "11" & x"3ca" => data <= x"f5";
            when "11" & x"3cb" => data <= x"00";
            when "11" & x"3cc" => data <= x"a2";
            when "11" & x"3cd" => data <= x"a0";
            when "11" & x"3ce" => data <= x"b1";
            when "11" & x"3cf" => data <= x"f2";
            when "11" & x"3d0" => data <= x"c9";
            when "11" & x"3d1" => data <= x"0d";
            when "11" & x"3d2" => data <= x"d0";
            when "11" & x"3d3" => data <= x"16";
            when "11" & x"3d4" => data <= x"98";
            when "11" & x"3d5" => data <= x"e8";
            when "11" & x"3d6" => data <= x"a0";
            when "11" & x"3d7" => data <= x"02";
            when "11" & x"3d8" => data <= x"20";
            when "11" & x"3d9" => data <= x"cb";
            when "11" & x"3da" => data <= x"99";
            when "11" & x"3db" => data <= x"20";
            when "11" & x"3dc" => data <= x"44";
            when "11" & x"3dd" => data <= x"b6";
            when "11" & x"3de" => data <= x"20";
            when "11" & x"3df" => data <= x"20";
            when "11" & x"3e0" => data <= x"44";
            when "11" & x"3e1" => data <= x"55";
            when "11" & x"3e2" => data <= x"54";
            when "11" & x"3e3" => data <= x"49";
            when "11" & x"3e4" => data <= x"4c";
            when "11" & x"3e5" => data <= x"53";
            when "11" & x"3e6" => data <= x"00";
            when "11" & x"3e7" => data <= x"4c";
            when "11" & x"3e8" => data <= x"e7";
            when "11" & x"3e9" => data <= x"ff";
            when "11" & x"3ea" => data <= x"98";
            when "11" & x"3eb" => data <= x"48";
            when "11" & x"3ec" => data <= x"20";
            when "11" & x"3ed" => data <= x"71";
            when "11" & x"3ee" => data <= x"86";
            when "11" & x"3ef" => data <= x"68";
            when "11" & x"3f0" => data <= x"a8";
            when "11" & x"3f1" => data <= x"a2";
            when "11" & x"3f2" => data <= x"92";
            when "11" & x"3f3" => data <= x"4c";
            when "11" & x"3f4" => data <= x"6e";
            when "11" & x"3f5" => data <= x"b4";
            when "11" & x"3f6" => data <= x"c8";
            when "11" & x"3f7" => data <= x"b1";
            when "11" & x"3f8" => data <= x"f2";
            when "11" & x"3f9" => data <= x"c9";
            when "11" & x"3fa" => data <= x"0d";
            when "11" & x"3fb" => data <= x"f0";
            when "11" & x"3fc" => data <= x"06";
            when "11" & x"3fd" => data <= x"c9";
            when "11" & x"3fe" => data <= x"20";
            when "11" & x"3ff" => data <= x"f0";
            when "11" & x"400" => data <= x"f0";
            when "11" & x"401" => data <= x"d0";
            when "11" & x"402" => data <= x"f3";
            when "11" & x"403" => data <= x"60";
            when "11" & x"404" => data <= x"20";
            when "11" & x"405" => data <= x"e7";
            when "11" & x"406" => data <= x"ff";
            when "11" & x"407" => data <= x"20";
            when "11" & x"408" => data <= x"44";
            when "11" & x"409" => data <= x"b6";
            when "11" & x"40a" => data <= x"53";
            when "11" & x"40b" => data <= x"50";
            when "11" & x"40c" => data <= x"49";
            when "11" & x"40d" => data <= x"20";
            when "11" & x"40e" => data <= x"30";
            when "11" & x"40f" => data <= x"2e";
            when "11" & x"410" => data <= x"30";
            when "11" & x"411" => data <= x"31";
            when "11" & x"412" => data <= x"00";
            when "11" & x"413" => data <= x"20";
            when "11" & x"414" => data <= x"e7";
            when "11" & x"415" => data <= x"ff";
            when "11" & x"416" => data <= x"a2";
            when "11" & x"417" => data <= x"00";
            when "11" & x"418" => data <= x"a9";
            when "11" & x"419" => data <= x"11";
            when "11" & x"41a" => data <= x"86";
            when "11" & x"41b" => data <= x"b5";
            when "11" & x"41c" => data <= x"85";
            when "11" & x"41d" => data <= x"bf";
            when "11" & x"41e" => data <= x"a2";
            when "11" & x"41f" => data <= x"00";
            when "11" & x"420" => data <= x"a9";
            when "11" & x"421" => data <= x"20";
            when "11" & x"422" => data <= x"20";
            when "11" & x"423" => data <= x"ee";
            when "11" & x"424" => data <= x"ff";
            when "11" & x"425" => data <= x"20";
            when "11" & x"426" => data <= x"ee";
            when "11" & x"427" => data <= x"ff";
            when "11" & x"428" => data <= x"20";
            when "11" & x"429" => data <= x"08";
            when "11" & x"42a" => data <= x"b7";
            when "11" & x"42b" => data <= x"20";
            when "11" & x"42c" => data <= x"e7";
            when "11" & x"42d" => data <= x"ff";
            when "11" & x"42e" => data <= x"c6";
            when "11" & x"42f" => data <= x"bf";
            when "11" & x"430" => data <= x"d0";
            when "11" & x"431" => data <= x"ee";
            when "11" & x"432" => data <= x"60";
            when "11" & x"433" => data <= x"20";
            when "11" & x"434" => data <= x"44";
            when "11" & x"435" => data <= x"b6";
            when "11" & x"436" => data <= x"44";
            when "11" & x"437" => data <= x"55";
            when "11" & x"438" => data <= x"54";
            when "11" & x"439" => data <= x"49";
            when "11" & x"43a" => data <= x"4c";
            when "11" & x"43b" => data <= x"53";
            when "11" & x"43c" => data <= x"20";
            when "11" & x"43d" => data <= x"62";
            when "11" & x"43e" => data <= x"79";
            when "11" & x"43f" => data <= x"20";
            when "11" & x"440" => data <= x"4d";
            when "11" & x"441" => data <= x"61";
            when "11" & x"442" => data <= x"72";
            when "11" & x"443" => data <= x"74";
            when "11" & x"444" => data <= x"69";
            when "11" & x"445" => data <= x"6e";
            when "11" & x"446" => data <= x"20";
            when "11" & x"447" => data <= x"4d";
            when "11" & x"448" => data <= x"61";
            when "11" & x"449" => data <= x"74";
            when "11" & x"44a" => data <= x"68";
            when "11" & x"44b" => data <= x"65";
            when "11" & x"44c" => data <= x"72";
            when "11" & x"44d" => data <= x"20";
            when "11" & x"44e" => data <= x"0a";
            when "11" & x"44f" => data <= x"0d";
            when "11" & x"450" => data <= x"4d";
            when "11" & x"451" => data <= x"4f";
            when "11" & x"452" => data <= x"44";
            when "11" & x"453" => data <= x"49";
            when "11" & x"454" => data <= x"46";
            when "11" & x"455" => data <= x"49";
            when "11" & x"456" => data <= x"45";
            when "11" & x"457" => data <= x"44";
            when "11" & x"458" => data <= x"20";
            when "11" & x"459" => data <= x"62";
            when "11" & x"45a" => data <= x"79";
            when "11" & x"45b" => data <= x"20";
            when "11" & x"45c" => data <= x"64";
            when "11" & x"45d" => data <= x"75";
            when "11" & x"45e" => data <= x"69";
            when "11" & x"45f" => data <= x"6b";
            when "11" & x"460" => data <= x"6b";
            when "11" & x"461" => data <= x"69";
            when "11" & x"462" => data <= x"65";
            when "11" & x"463" => data <= x"20";
            when "11" & x"464" => data <= x"32";
            when "11" & x"465" => data <= x"30";
            when "11" & x"466" => data <= x"31";
            when "11" & x"467" => data <= x"35";
            when "11" & x"468" => data <= x"00";
            when "11" & x"469" => data <= x"4c";
            when "11" & x"46a" => data <= x"e7";
            when "11" & x"46b" => data <= x"ff";
            when "11" & x"46c" => data <= x"a2";
            when "11" & x"46d" => data <= x"fd";
            when "11" & x"46e" => data <= x"98";
            when "11" & x"46f" => data <= x"48";
            when "11" & x"470" => data <= x"e8";
            when "11" & x"471" => data <= x"e8";
            when "11" & x"472" => data <= x"68";
            when "11" & x"473" => data <= x"48";
            when "11" & x"474" => data <= x"a8";
            when "11" & x"475" => data <= x"20";
            when "11" & x"476" => data <= x"b0";
            when "11" & x"477" => data <= x"b4";
            when "11" & x"478" => data <= x"e8";
            when "11" & x"479" => data <= x"bd";
            when "11" & x"47a" => data <= x"2b";
            when "11" & x"47b" => data <= x"b3";
            when "11" & x"47c" => data <= x"30";
            when "11" & x"47d" => data <= x"28";
            when "11" & x"47e" => data <= x"86";
            when "11" & x"47f" => data <= x"b5";
            when "11" & x"480" => data <= x"ca";
            when "11" & x"481" => data <= x"88";
            when "11" & x"482" => data <= x"e8";
            when "11" & x"483" => data <= x"c8";
            when "11" & x"484" => data <= x"bd";
            when "11" & x"485" => data <= x"2b";
            when "11" & x"486" => data <= x"b3";
            when "11" & x"487" => data <= x"30";
            when "11" & x"488" => data <= x"16";
            when "11" & x"489" => data <= x"51";
            when "11" & x"48a" => data <= x"f2";
            when "11" & x"48b" => data <= x"29";
            when "11" & x"48c" => data <= x"5f";
            when "11" & x"48d" => data <= x"f0";
            when "11" & x"48e" => data <= x"f3";
            when "11" & x"48f" => data <= x"ca";
            when "11" & x"490" => data <= x"e8";
            when "11" & x"491" => data <= x"bd";
            when "11" & x"492" => data <= x"2b";
            when "11" & x"493" => data <= x"b3";
            when "11" & x"494" => data <= x"10";
            when "11" & x"495" => data <= x"fa";
            when "11" & x"496" => data <= x"b1";
            when "11" & x"497" => data <= x"f2";
            when "11" & x"498" => data <= x"c9";
            when "11" & x"499" => data <= x"2e";
            when "11" & x"49a" => data <= x"d0";
            when "11" & x"49b" => data <= x"d4";
            when "11" & x"49c" => data <= x"c8";
            when "11" & x"49d" => data <= x"b0";
            when "11" & x"49e" => data <= x"07";
            when "11" & x"49f" => data <= x"b1";
            when "11" & x"4a0" => data <= x"f2";
            when "11" & x"4a1" => data <= x"20";
            when "11" & x"4a2" => data <= x"ee";
            when "11" & x"4a3" => data <= x"82";
            when "11" & x"4a4" => data <= x"90";
            when "11" & x"4a5" => data <= x"ca";
            when "11" & x"4a6" => data <= x"68";
            when "11" & x"4a7" => data <= x"bd";
            when "11" & x"4a8" => data <= x"2b";
            when "11" & x"4a9" => data <= x"b3";
            when "11" & x"4aa" => data <= x"48";
            when "11" & x"4ab" => data <= x"bd";
            when "11" & x"4ac" => data <= x"2c";
            when "11" & x"4ad" => data <= x"b3";
            when "11" & x"4ae" => data <= x"48";
            when "11" & x"4af" => data <= x"60";
            when "11" & x"4b0" => data <= x"b1";
            when "11" & x"4b1" => data <= x"f2";
            when "11" & x"4b2" => data <= x"c9";
            when "11" & x"4b3" => data <= x"0d";
            when "11" & x"4b4" => data <= x"f0";
            when "11" & x"4b5" => data <= x"08";
            when "11" & x"4b6" => data <= x"c8";
            when "11" & x"4b7" => data <= x"f0";
            when "11" & x"4b8" => data <= x"07";
            when "11" & x"4b9" => data <= x"c9";
            when "11" & x"4ba" => data <= x"20";
            when "11" & x"4bb" => data <= x"f0";
            when "11" & x"4bc" => data <= x"f3";
            when "11" & x"4bd" => data <= x"18";
            when "11" & x"4be" => data <= x"88";
            when "11" & x"4bf" => data <= x"60";
            when "11" & x"4c0" => data <= x"4c";
            when "11" & x"4c1" => data <= x"f5";
            when "11" & x"4c2" => data <= x"b6";
            when "11" & x"4c3" => data <= x"98";
            when "11" & x"4c4" => data <= x"48";
            when "11" & x"4c5" => data <= x"a9";
            when "11" & x"4c6" => data <= x"00";
            when "11" & x"4c7" => data <= x"8d";
            when "11" & x"4c8" => data <= x"55";
            when "11" & x"4c9" => data <= x"0d";
            when "11" & x"4ca" => data <= x"8d";
            when "11" & x"4cb" => data <= x"56";
            when "11" & x"4cc" => data <= x"0d";
            when "11" & x"4cd" => data <= x"20";
            when "11" & x"4ce" => data <= x"b0";
            when "11" & x"4cf" => data <= x"b4";
            when "11" & x"4d0" => data <= x"b0";
            when "11" & x"4d1" => data <= x"62";
            when "11" & x"4d2" => data <= x"b1";
            when "11" & x"4d3" => data <= x"f2";
            when "11" & x"4d4" => data <= x"c9";
            when "11" & x"4d5" => data <= x"0d";
            when "11" & x"4d6" => data <= x"f0";
            when "11" & x"4d7" => data <= x"5c";
            when "11" & x"4d8" => data <= x"38";
            when "11" & x"4d9" => data <= x"e9";
            when "11" & x"4da" => data <= x"30";
            when "11" & x"4db" => data <= x"30";
            when "11" & x"4dc" => data <= x"57";
            when "11" & x"4dd" => data <= x"c9";
            when "11" & x"4de" => data <= x"0a";
            when "11" & x"4df" => data <= x"b0";
            when "11" & x"4e0" => data <= x"53";
            when "11" & x"4e1" => data <= x"48";
            when "11" & x"4e2" => data <= x"ad";
            when "11" & x"4e3" => data <= x"55";
            when "11" & x"4e4" => data <= x"0d";
            when "11" & x"4e5" => data <= x"0a";
            when "11" & x"4e6" => data <= x"48";
            when "11" & x"4e7" => data <= x"2e";
            when "11" & x"4e8" => data <= x"56";
            when "11" & x"4e9" => data <= x"0d";
            when "11" & x"4ea" => data <= x"ae";
            when "11" & x"4eb" => data <= x"56";
            when "11" & x"4ec" => data <= x"0d";
            when "11" & x"4ed" => data <= x"0a";
            when "11" & x"4ee" => data <= x"2e";
            when "11" & x"4ef" => data <= x"56";
            when "11" & x"4f0" => data <= x"0d";
            when "11" & x"4f1" => data <= x"0a";
            when "11" & x"4f2" => data <= x"2e";
            when "11" & x"4f3" => data <= x"56";
            when "11" & x"4f4" => data <= x"0d";
            when "11" & x"4f5" => data <= x"8d";
            when "11" & x"4f6" => data <= x"55";
            when "11" & x"4f7" => data <= x"0d";
            when "11" & x"4f8" => data <= x"68";
            when "11" & x"4f9" => data <= x"6d";
            when "11" & x"4fa" => data <= x"55";
            when "11" & x"4fb" => data <= x"0d";
            when "11" & x"4fc" => data <= x"8d";
            when "11" & x"4fd" => data <= x"55";
            when "11" & x"4fe" => data <= x"0d";
            when "11" & x"4ff" => data <= x"8a";
            when "11" & x"500" => data <= x"6d";
            when "11" & x"501" => data <= x"56";
            when "11" & x"502" => data <= x"0d";
            when "11" & x"503" => data <= x"aa";
            when "11" & x"504" => data <= x"68";
            when "11" & x"505" => data <= x"6d";
            when "11" & x"506" => data <= x"55";
            when "11" & x"507" => data <= x"0d";
            when "11" & x"508" => data <= x"8d";
            when "11" & x"509" => data <= x"55";
            when "11" & x"50a" => data <= x"0d";
            when "11" & x"50b" => data <= x"8a";
            when "11" & x"50c" => data <= x"69";
            when "11" & x"50d" => data <= x"00";
            when "11" & x"50e" => data <= x"8d";
            when "11" & x"50f" => data <= x"56";
            when "11" & x"510" => data <= x"0d";
            when "11" & x"511" => data <= x"c9";
            when "11" & x"512" => data <= x"02";
            when "11" & x"513" => data <= x"b0";
            when "11" & x"514" => data <= x"1f";
            when "11" & x"515" => data <= x"c8";
            when "11" & x"516" => data <= x"f0";
            when "11" & x"517" => data <= x"1c";
            when "11" & x"518" => data <= x"b1";
            when "11" & x"519" => data <= x"f2";
            when "11" & x"51a" => data <= x"c9";
            when "11" & x"51b" => data <= x"0d";
            when "11" & x"51c" => data <= x"f0";
            when "11" & x"51d" => data <= x"04";
            when "11" & x"51e" => data <= x"c9";
            when "11" & x"51f" => data <= x"20";
            when "11" & x"520" => data <= x"d0";
            when "11" & x"521" => data <= x"b6";
            when "11" & x"522" => data <= x"ae";
            when "11" & x"523" => data <= x"55";
            when "11" & x"524" => data <= x"0d";
            when "11" & x"525" => data <= x"ad";
            when "11" & x"526" => data <= x"56";
            when "11" & x"527" => data <= x"0d";
            when "11" & x"528" => data <= x"f0";
            when "11" & x"529" => data <= x"04";
            when "11" & x"52a" => data <= x"e8";
            when "11" & x"52b" => data <= x"f0";
            when "11" & x"52c" => data <= x"07";
            when "11" & x"52d" => data <= x"ca";
            when "11" & x"52e" => data <= x"68";
            when "11" & x"52f" => data <= x"ad";
            when "11" & x"530" => data <= x"56";
            when "11" & x"531" => data <= x"0d";
            when "11" & x"532" => data <= x"18";
            when "11" & x"533" => data <= x"60";
            when "11" & x"534" => data <= x"68";
            when "11" & x"535" => data <= x"a8";
            when "11" & x"536" => data <= x"a9";
            when "11" & x"537" => data <= x"00";
            when "11" & x"538" => data <= x"aa";
            when "11" & x"539" => data <= x"38";
            when "11" & x"53a" => data <= x"60";
            when "11" & x"53b" => data <= x"a9";
            when "11" & x"53c" => data <= x"0d";
            when "11" & x"53d" => data <= x"8d";
            when "11" & x"53e" => data <= x"5d";
            when "11" & x"53f" => data <= x"0d";
            when "11" & x"540" => data <= x"a2";
            when "11" & x"541" => data <= x"00";
            when "11" & x"542" => data <= x"8e";
            when "11" & x"543" => data <= x"5e";
            when "11" & x"544" => data <= x"0d";
            when "11" & x"545" => data <= x"20";
            when "11" & x"546" => data <= x"b0";
            when "11" & x"547" => data <= x"b4";
            when "11" & x"548" => data <= x"b0";
            when "11" & x"549" => data <= x"49";
            when "11" & x"54a" => data <= x"c9";
            when "11" & x"54b" => data <= x"22";
            when "11" & x"54c" => data <= x"d0";
            when "11" & x"54d" => data <= x"04";
            when "11" & x"54e" => data <= x"c8";
            when "11" & x"54f" => data <= x"8d";
            when "11" & x"550" => data <= x"5d";
            when "11" & x"551" => data <= x"0d";
            when "11" & x"552" => data <= x"b1";
            when "11" & x"553" => data <= x"f2";
            when "11" & x"554" => data <= x"c9";
            when "11" & x"555" => data <= x"0d";
            when "11" & x"556" => data <= x"f0";
            when "11" & x"557" => data <= x"2c";
            when "11" & x"558" => data <= x"c9";
            when "11" & x"559" => data <= x"20";
            when "11" & x"55a" => data <= x"d0";
            when "11" & x"55b" => data <= x"0b";
            when "11" & x"55c" => data <= x"90";
            when "11" & x"55d" => data <= x"52";
            when "11" & x"55e" => data <= x"ad";
            when "11" & x"55f" => data <= x"5d";
            when "11" & x"560" => data <= x"0d";
            when "11" & x"561" => data <= x"c9";
            when "11" & x"562" => data <= x"22";
            when "11" & x"563" => data <= x"d0";
            when "11" & x"564" => data <= x"28";
            when "11" & x"565" => data <= x"a9";
            when "11" & x"566" => data <= x"20";
            when "11" & x"567" => data <= x"c9";
            when "11" & x"568" => data <= x"22";
            when "11" & x"569" => data <= x"f0";
            when "11" & x"56a" => data <= x"19";
            when "11" & x"56b" => data <= x"c9";
            when "11" & x"56c" => data <= x"2a";
            when "11" & x"56d" => data <= x"f0";
            when "11" & x"56e" => data <= x"31";
            when "11" & x"56f" => data <= x"c9";
            when "11" & x"570" => data <= x"61";
            when "11" & x"571" => data <= x"90";
            when "11" & x"572" => data <= x"06";
            when "11" & x"573" => data <= x"c9";
            when "11" & x"574" => data <= x"7b";
            when "11" & x"575" => data <= x"b0";
            when "11" & x"576" => data <= x"02";
            when "11" & x"577" => data <= x"49";
            when "11" & x"578" => data <= x"20";
            when "11" & x"579" => data <= x"9d";
            when "11" & x"57a" => data <= x"5f";
            when "11" & x"57b" => data <= x"0d";
            when "11" & x"57c" => data <= x"c8";
            when "11" & x"57d" => data <= x"e8";
            when "11" & x"57e" => data <= x"e0";
            when "11" & x"57f" => data <= x"0c";
            when "11" & x"580" => data <= x"d0";
            when "11" & x"581" => data <= x"d0";
            when "11" & x"582" => data <= x"b1";
            when "11" & x"583" => data <= x"f2";
            when "11" & x"584" => data <= x"cd";
            when "11" & x"585" => data <= x"5d";
            when "11" & x"586" => data <= x"0d";
            when "11" & x"587" => data <= x"d0";
            when "11" & x"588" => data <= x"27";
            when "11" & x"589" => data <= x"c9";
            when "11" & x"58a" => data <= x"0d";
            when "11" & x"58b" => data <= x"f0";
            when "11" & x"58c" => data <= x"06";
            when "11" & x"58d" => data <= x"c8";
            when "11" & x"58e" => data <= x"20";
            when "11" & x"58f" => data <= x"b0";
            when "11" & x"590" => data <= x"b4";
            when "11" & x"591" => data <= x"90";
            when "11" & x"592" => data <= x"1d";
            when "11" & x"593" => data <= x"8e";
            when "11" & x"594" => data <= x"5c";
            when "11" & x"595" => data <= x"0d";
            when "11" & x"596" => data <= x"e0";
            when "11" & x"597" => data <= x"0c";
            when "11" & x"598" => data <= x"f0";
            when "11" & x"599" => data <= x"05";
            when "11" & x"59a" => data <= x"a9";
            when "11" & x"59b" => data <= x"00";
            when "11" & x"59c" => data <= x"9d";
            when "11" & x"59d" => data <= x"5f";
            when "11" & x"59e" => data <= x"0d";
            when "11" & x"59f" => data <= x"60";
            when "11" & x"5a0" => data <= x"8d";
            when "11" & x"5a1" => data <= x"5e";
            when "11" & x"5a2" => data <= x"0d";
            when "11" & x"5a3" => data <= x"ad";
            when "11" & x"5a4" => data <= x"5d";
            when "11" & x"5a5" => data <= x"0d";
            when "11" & x"5a6" => data <= x"c9";
            when "11" & x"5a7" => data <= x"0d";
            when "11" & x"5a8" => data <= x"f0";
            when "11" & x"5a9" => data <= x"e3";
            when "11" & x"5aa" => data <= x"c8";
            when "11" & x"5ab" => data <= x"b1";
            when "11" & x"5ac" => data <= x"f2";
            when "11" & x"5ad" => data <= x"4c";
            when "11" & x"5ae" => data <= x"84";
            when "11" & x"5af" => data <= x"b5";
            when "11" & x"5b0" => data <= x"4c";
            when "11" & x"5b1" => data <= x"f5";
            when "11" & x"5b2" => data <= x"b6";
            when "11" & x"5b3" => data <= x"a0";
            when "11" & x"5b4" => data <= x"00";
            when "11" & x"5b5" => data <= x"ae";
            when "11" & x"5b6" => data <= x"5c";
            when "11" & x"5b7" => data <= x"0d";
            when "11" & x"5b8" => data <= x"f0";
            when "11" & x"5b9" => data <= x"17";
            when "11" & x"5ba" => data <= x"b1";
            when "11" & x"5bb" => data <= x"f2";
            when "11" & x"5bc" => data <= x"f0";
            when "11" & x"5bd" => data <= x"25";
            when "11" & x"5be" => data <= x"c9";
            when "11" & x"5bf" => data <= x"61";
            when "11" & x"5c0" => data <= x"90";
            when "11" & x"5c1" => data <= x"06";
            when "11" & x"5c2" => data <= x"c9";
            when "11" & x"5c3" => data <= x"7b";
            when "11" & x"5c4" => data <= x"b0";
            when "11" & x"5c5" => data <= x"02";
            when "11" & x"5c6" => data <= x"49";
            when "11" & x"5c7" => data <= x"20";
            when "11" & x"5c8" => data <= x"d9";
            when "11" & x"5c9" => data <= x"5f";
            when "11" & x"5ca" => data <= x"0d";
            when "11" & x"5cb" => data <= x"d0";
            when "11" & x"5cc" => data <= x"16";
            when "11" & x"5cd" => data <= x"c8";
            when "11" & x"5ce" => data <= x"ca";
            when "11" & x"5cf" => data <= x"d0";
            when "11" & x"5d0" => data <= x"e9";
            when "11" & x"5d1" => data <= x"b1";
            when "11" & x"5d2" => data <= x"f2";
            when "11" & x"5d3" => data <= x"f0";
            when "11" & x"5d4" => data <= x"0c";
            when "11" & x"5d5" => data <= x"ad";
            when "11" & x"5d6" => data <= x"5c";
            when "11" & x"5d7" => data <= x"0d";
            when "11" & x"5d8" => data <= x"c9";
            when "11" & x"5d9" => data <= x"0c";
            when "11" & x"5da" => data <= x"f0";
            when "11" & x"5db" => data <= x"05";
            when "11" & x"5dc" => data <= x"ad";
            when "11" & x"5dd" => data <= x"5e";
            when "11" & x"5de" => data <= x"0d";
            when "11" & x"5df" => data <= x"f0";
            when "11" & x"5e0" => data <= x"02";
            when "11" & x"5e1" => data <= x"18";
            when "11" & x"5e2" => data <= x"60";
            when "11" & x"5e3" => data <= x"38";
            when "11" & x"5e4" => data <= x"60";
            when "11" & x"5e5" => data <= x"b0";
            when "11" & x"5e6" => data <= x"05";
            when "11" & x"5e7" => data <= x"a9";
            when "11" & x"5e8" => data <= x"20";
            when "11" & x"5e9" => data <= x"20";
            when "11" & x"5ea" => data <= x"ee";
            when "11" & x"5eb" => data <= x"ff";
            when "11" & x"5ec" => data <= x"a2";
            when "11" & x"5ed" => data <= x"20";
            when "11" & x"5ee" => data <= x"a0";
            when "11" & x"5ef" => data <= x"04";
            when "11" & x"5f0" => data <= x"ad";
            when "11" & x"5f1" => data <= x"56";
            when "11" & x"5f2" => data <= x"0d";
            when "11" & x"5f3" => data <= x"20";
            when "11" & x"5f4" => data <= x"26";
            when "11" & x"5f5" => data <= x"b6";
            when "11" & x"5f6" => data <= x"ad";
            when "11" & x"5f7" => data <= x"55";
            when "11" & x"5f8" => data <= x"0d";
            when "11" & x"5f9" => data <= x"20";
            when "11" & x"5fa" => data <= x"26";
            when "11" & x"5fb" => data <= x"b6";
            when "11" & x"5fc" => data <= x"a9";
            when "11" & x"5fd" => data <= x"20";
            when "11" & x"5fe" => data <= x"20";
            when "11" & x"5ff" => data <= x"ee";
            when "11" & x"600" => data <= x"ff";
            when "11" & x"601" => data <= x"a0";
            when "11" & x"602" => data <= x"00";
            when "11" & x"603" => data <= x"b1";
            when "11" & x"604" => data <= x"f2";
            when "11" & x"605" => data <= x"f0";
            when "11" & x"606" => data <= x"08";
            when "11" & x"607" => data <= x"20";
            when "11" & x"608" => data <= x"ee";
            when "11" & x"609" => data <= x"ff";
            when "11" & x"60a" => data <= x"c8";
            when "11" & x"60b" => data <= x"c0";
            when "11" & x"60c" => data <= x"0c";
            when "11" & x"60d" => data <= x"d0";
            when "11" & x"60e" => data <= x"f4";
            when "11" & x"60f" => data <= x"a9";
            when "11" & x"610" => data <= x"20";
            when "11" & x"611" => data <= x"20";
            when "11" & x"612" => data <= x"ee";
            when "11" & x"613" => data <= x"ff";
            when "11" & x"614" => data <= x"c8";
            when "11" & x"615" => data <= x"c0";
            when "11" & x"616" => data <= x"0d";
            when "11" & x"617" => data <= x"d0";
            when "11" & x"618" => data <= x"f8";
            when "11" & x"619" => data <= x"aa";
            when "11" & x"61a" => data <= x"a0";
            when "11" & x"61b" => data <= x"0f";
            when "11" & x"61c" => data <= x"b1";
            when "11" & x"61d" => data <= x"f2";
            when "11" & x"61e" => data <= x"d0";
            when "11" & x"61f" => data <= x"02";
            when "11" & x"620" => data <= x"a2";
            when "11" & x"621" => data <= x"50";
            when "11" & x"622" => data <= x"8a";
            when "11" & x"623" => data <= x"4c";
            when "11" & x"624" => data <= x"ee";
            when "11" & x"625" => data <= x"ff";
            when "11" & x"626" => data <= x"48";
            when "11" & x"627" => data <= x"4a";
            when "11" & x"628" => data <= x"4a";
            when "11" & x"629" => data <= x"4a";
            when "11" & x"62a" => data <= x"4a";
            when "11" & x"62b" => data <= x"20";
            when "11" & x"62c" => data <= x"2f";
            when "11" & x"62d" => data <= x"b6";
            when "11" & x"62e" => data <= x"68";
            when "11" & x"62f" => data <= x"29";
            when "11" & x"630" => data <= x"0f";
            when "11" & x"631" => data <= x"f0";
            when "11" & x"632" => data <= x"08";
            when "11" & x"633" => data <= x"a2";
            when "11" & x"634" => data <= x"30";
            when "11" & x"635" => data <= x"18";
            when "11" & x"636" => data <= x"69";
            when "11" & x"637" => data <= x"30";
            when "11" & x"638" => data <= x"4c";
            when "11" & x"639" => data <= x"ee";
            when "11" & x"63a" => data <= x"ff";
            when "11" & x"63b" => data <= x"88";
            when "11" & x"63c" => data <= x"d0";
            when "11" & x"63d" => data <= x"02";
            when "11" & x"63e" => data <= x"a2";
            when "11" & x"63f" => data <= x"30";
            when "11" & x"640" => data <= x"8a";
            when "11" & x"641" => data <= x"4c";
            when "11" & x"642" => data <= x"ee";
            when "11" & x"643" => data <= x"ff";
            when "11" & x"644" => data <= x"a2";
            when "11" & x"645" => data <= x"00";
            when "11" & x"646" => data <= x"68";
            when "11" & x"647" => data <= x"85";
            when "11" & x"648" => data <= x"a0";
            when "11" & x"649" => data <= x"68";
            when "11" & x"64a" => data <= x"85";
            when "11" & x"64b" => data <= x"a1";
            when "11" & x"64c" => data <= x"a0";
            when "11" & x"64d" => data <= x"00";
            when "11" & x"64e" => data <= x"f0";
            when "11" & x"64f" => data <= x"07";
            when "11" & x"650" => data <= x"b1";
            when "11" & x"651" => data <= x"a0";
            when "11" & x"652" => data <= x"f0";
            when "11" & x"653" => data <= x"0b";
            when "11" & x"654" => data <= x"20";
            when "11" & x"655" => data <= x"66";
            when "11" & x"656" => data <= x"b6";
            when "11" & x"657" => data <= x"e6";
            when "11" & x"658" => data <= x"a0";
            when "11" & x"659" => data <= x"d0";
            when "11" & x"65a" => data <= x"f5";
            when "11" & x"65b" => data <= x"e6";
            when "11" & x"65c" => data <= x"a1";
            when "11" & x"65d" => data <= x"d0";
            when "11" & x"65e" => data <= x"f1";
            when "11" & x"65f" => data <= x"a5";
            when "11" & x"660" => data <= x"a1";
            when "11" & x"661" => data <= x"48";
            when "11" & x"662" => data <= x"a5";
            when "11" & x"663" => data <= x"a0";
            when "11" & x"664" => data <= x"48";
            when "11" & x"665" => data <= x"60";
            when "11" & x"666" => data <= x"e0";
            when "11" & x"667" => data <= x"00";
            when "11" & x"668" => data <= x"d0";
            when "11" & x"669" => data <= x"03";
            when "11" & x"66a" => data <= x"4c";
            when "11" & x"66b" => data <= x"ee";
            when "11" & x"66c" => data <= x"ff";
            when "11" & x"66d" => data <= x"9d";
            when "11" & x"66e" => data <= x"00";
            when "11" & x"66f" => data <= x"01";
            when "11" & x"670" => data <= x"e8";
            when "11" & x"671" => data <= x"60";
            when "11" & x"672" => data <= x"08";
            when "11" & x"673" => data <= x"10";
            when "11" & x"674" => data <= x"1c";
            when "11" & x"675" => data <= x"22";
            when "11" & x"676" => data <= x"43";
            when "11" & x"677" => data <= x"49";
            when "11" & x"678" => data <= x"4f";
            when "11" & x"679" => data <= x"58";
            when "11" & x"67a" => data <= x"28";
            when "11" & x"67b" => data <= x"3c";
            when "11" & x"67c" => data <= x"64";
            when "11" & x"67d" => data <= x"72";
            when "11" & x"67e" => data <= x"76";
            when "11" & x"67f" => data <= x"3e";
            when "11" & x"680" => data <= x"29";
            when "11" & x"681" => data <= x"00";
            when "11" & x"682" => data <= x"3c";
            when "11" & x"683" => data <= x"64";
            when "11" & x"684" => data <= x"6e";
            when "11" & x"685" => data <= x"6f";
            when "11" & x"686" => data <= x"3e";
            when "11" & x"687" => data <= x"2f";
            when "11" & x"688" => data <= x"3c";
            when "11" & x"689" => data <= x"64";
            when "11" & x"68a" => data <= x"73";
            when "11" & x"68b" => data <= x"70";
            when "11" & x"68c" => data <= x"3e";
            when "11" & x"68d" => data <= x"00";
            when "11" & x"68e" => data <= x"3c";
            when "11" & x"68f" => data <= x"64";
            when "11" & x"690" => data <= x"6e";
            when "11" & x"691" => data <= x"6f";
            when "11" & x"692" => data <= x"3e";
            when "11" & x"693" => data <= x"00";
            when "11" & x"694" => data <= x"28";
            when "11" & x"695" => data <= x"28";
            when "11" & x"696" => data <= x"3c";
            when "11" & x"697" => data <= x"66";
            when "11" & x"698" => data <= x"72";
            when "11" & x"699" => data <= x"6f";
            when "11" & x"69a" => data <= x"6d";
            when "11" & x"69b" => data <= x"20";
            when "11" & x"69c" => data <= x"64";
            when "11" & x"69d" => data <= x"6e";
            when "11" & x"69e" => data <= x"6f";
            when "11" & x"69f" => data <= x"3e";
            when "11" & x"6a0" => data <= x"29";
            when "11" & x"6a1" => data <= x"20";
            when "11" & x"6a2" => data <= x"3c";
            when "11" & x"6a3" => data <= x"74";
            when "11" & x"6a4" => data <= x"6f";
            when "11" & x"6a5" => data <= x"20";
            when "11" & x"6a6" => data <= x"64";
            when "11" & x"6a7" => data <= x"6e";
            when "11" & x"6a8" => data <= x"6f";
            when "11" & x"6a9" => data <= x"3e";
            when "11" & x"6aa" => data <= x"29";
            when "11" & x"6ab" => data <= x"20";
            when "11" & x"6ac" => data <= x"28";
            when "11" & x"6ad" => data <= x"3c";
            when "11" & x"6ae" => data <= x"61";
            when "11" & x"6af" => data <= x"64";
            when "11" & x"6b0" => data <= x"73";
            when "11" & x"6b1" => data <= x"70";
            when "11" & x"6b2" => data <= x"3e";
            when "11" & x"6b3" => data <= x"29";
            when "11" & x"6b4" => data <= x"00";
            when "11" & x"6b5" => data <= x"3c";
            when "11" & x"6b6" => data <= x"64";
            when "11" & x"6b7" => data <= x"72";
            when "11" & x"6b8" => data <= x"76";
            when "11" & x"6b9" => data <= x"3e";
            when "11" & x"6ba" => data <= x"00";
            when "11" & x"6bb" => data <= x"3c";
            when "11" & x"6bc" => data <= x"66";
            when "11" & x"6bd" => data <= x"73";
            when "11" & x"6be" => data <= x"70";
            when "11" & x"6bf" => data <= x"3e";
            when "11" & x"6c0" => data <= x"00";
            when "11" & x"6c1" => data <= x"28";
            when "11" & x"6c2" => data <= x"3c";
            when "11" & x"6c3" => data <= x"6d";
            when "11" & x"6c4" => data <= x"6f";
            when "11" & x"6c5" => data <= x"64";
            when "11" & x"6c6" => data <= x"65";
            when "11" & x"6c7" => data <= x"3e";
            when "11" & x"6c8" => data <= x"29";
            when "11" & x"6c9" => data <= x"00";
            when "11" & x"6ca" => data <= x"28";
            when "11" & x"6cb" => data <= x"3c";
            when "11" & x"6cc" => data <= x"72";
            when "11" & x"6cd" => data <= x"6f";
            when "11" & x"6ce" => data <= x"6d";
            when "11" & x"6cf" => data <= x"3e";
            when "11" & x"6d0" => data <= x"29";
            when "11" & x"6d1" => data <= x"00";
            when "11" & x"6d2" => data <= x"48";
            when "11" & x"6d3" => data <= x"4a";
            when "11" & x"6d4" => data <= x"4a";
            when "11" & x"6d5" => data <= x"4a";
            when "11" & x"6d6" => data <= x"4a";
            when "11" & x"6d7" => data <= x"20";
            when "11" & x"6d8" => data <= x"dd";
            when "11" & x"6d9" => data <= x"b6";
            when "11" & x"6da" => data <= x"68";
            when "11" & x"6db" => data <= x"29";
            when "11" & x"6dc" => data <= x"0f";
            when "11" & x"6dd" => data <= x"a8";
            when "11" & x"6de" => data <= x"f0";
            when "11" & x"6df" => data <= x"14";
            when "11" & x"6e0" => data <= x"a9";
            when "11" & x"6e1" => data <= x"20";
            when "11" & x"6e2" => data <= x"20";
            when "11" & x"6e3" => data <= x"66";
            when "11" & x"6e4" => data <= x"b6";
            when "11" & x"6e5" => data <= x"b9";
            when "11" & x"6e6" => data <= x"71";
            when "11" & x"6e7" => data <= x"b6";
            when "11" & x"6e8" => data <= x"a8";
            when "11" & x"6e9" => data <= x"b9";
            when "11" & x"6ea" => data <= x"72";
            when "11" & x"6eb" => data <= x"b6";
            when "11" & x"6ec" => data <= x"f0";
            when "11" & x"6ed" => data <= x"06";
            when "11" & x"6ee" => data <= x"20";
            when "11" & x"6ef" => data <= x"66";
            when "11" & x"6f0" => data <= x"b6";
            when "11" & x"6f1" => data <= x"c8";
            when "11" & x"6f2" => data <= x"d0";
            when "11" & x"6f3" => data <= x"f5";
            when "11" & x"6f4" => data <= x"60";
            when "11" & x"6f5" => data <= x"a2";
            when "11" & x"6f6" => data <= x"00";
            when "11" & x"6f7" => data <= x"8e";
            when "11" & x"6f8" => data <= x"00";
            when "11" & x"6f9" => data <= x"01";
            when "11" & x"6fa" => data <= x"e8";
            when "11" & x"6fb" => data <= x"20";
            when "11" & x"6fc" => data <= x"46";
            when "11" & x"6fd" => data <= x"b6";
            when "11" & x"6fe" => data <= x"1a";
            when "11" & x"6ff" => data <= x"53";
            when "11" & x"700" => data <= x"79";
            when "11" & x"701" => data <= x"6e";
            when "11" & x"702" => data <= x"74";
            when "11" & x"703" => data <= x"61";
            when "11" & x"704" => data <= x"78";
            when "11" & x"705" => data <= x"3a";
            when "11" & x"706" => data <= x"20";
            when "11" & x"707" => data <= x"00";
            when "11" & x"708" => data <= x"a4";
            when "11" & x"709" => data <= x"b5";
            when "11" & x"70a" => data <= x"b9";
            when "11" & x"70b" => data <= x"2b";
            when "11" & x"70c" => data <= x"b3";
            when "11" & x"70d" => data <= x"30";
            when "11" & x"70e" => data <= x"06";
            when "11" & x"70f" => data <= x"20";
            when "11" & x"710" => data <= x"66";
            when "11" & x"711" => data <= x"b6";
            when "11" & x"712" => data <= x"c8";
            when "11" & x"713" => data <= x"d0";
            when "11" & x"714" => data <= x"f5";
            when "11" & x"715" => data <= x"c8";
            when "11" & x"716" => data <= x"c8";
            when "11" & x"717" => data <= x"b9";
            when "11" & x"718" => data <= x"2b";
            when "11" & x"719" => data <= x"b3";
            when "11" & x"71a" => data <= x"c8";
            when "11" & x"71b" => data <= x"84";
            when "11" & x"71c" => data <= x"b5";
            when "11" & x"71d" => data <= x"20";
            when "11" & x"71e" => data <= x"d2";
            when "11" & x"71f" => data <= x"b6";
            when "11" & x"720" => data <= x"e0";
            when "11" & x"721" => data <= x"00";
            when "11" & x"722" => data <= x"f0";
            when "11" & x"723" => data <= x"08";
            when "11" & x"724" => data <= x"a9";
            when "11" & x"725" => data <= x"00";
            when "11" & x"726" => data <= x"9d";
            when "11" & x"727" => data <= x"00";
            when "11" & x"728" => data <= x"01";
            when "11" & x"729" => data <= x"4c";
            when "11" & x"72a" => data <= x"00";
            when "11" & x"72b" => data <= x"01";
            when "11" & x"72c" => data <= x"60";
            when "11" & x"72d" => data <= x"4c";
            when "11" & x"72e" => data <= x"f5";
            when "11" & x"72f" => data <= x"b6";
            when "11" & x"730" => data <= x"20";
            when "11" & x"731" => data <= x"b0";
            when "11" & x"732" => data <= x"b4";
            when "11" & x"733" => data <= x"b0";
            when "11" & x"734" => data <= x"17";
            when "11" & x"735" => data <= x"20";
            when "11" & x"736" => data <= x"c3";
            when "11" & x"737" => data <= x"b4";
            when "11" & x"738" => data <= x"b0";
            when "11" & x"739" => data <= x"bb";
            when "11" & x"73a" => data <= x"48";
            when "11" & x"73b" => data <= x"20";
            when "11" & x"73c" => data <= x"b0";
            when "11" & x"73d" => data <= x"b4";
            when "11" & x"73e" => data <= x"68";
            when "11" & x"73f" => data <= x"90";
            when "11" & x"740" => data <= x"b4";
            when "11" & x"741" => data <= x"d0";
            when "11" & x"742" => data <= x"26";
            when "11" & x"743" => data <= x"8a";
            when "11" & x"744" => data <= x"8d";
            when "11" & x"745" => data <= x"5b";
            when "11" & x"746" => data <= x"0d";
            when "11" & x"747" => data <= x"c9";
            when "11" & x"748" => data <= x"04";
            when "11" & x"749" => data <= x"b0";
            when "11" & x"74a" => data <= x"1e";
            when "11" & x"74b" => data <= x"60";
            when "11" & x"74c" => data <= x"a5";
            when "11" & x"74d" => data <= x"cf";
            when "11" & x"74e" => data <= x"60";
            when "11" & x"74f" => data <= x"20";
            when "11" & x"750" => data <= x"b0";
            when "11" & x"751" => data <= x"b4";
            when "11" & x"752" => data <= x"b0";
            when "11" & x"753" => data <= x"a1";
            when "11" & x"754" => data <= x"20";
            when "11" & x"755" => data <= x"c3";
            when "11" & x"756" => data <= x"b4";
            when "11" & x"757" => data <= x"b0";
            when "11" & x"758" => data <= x"9c";
            when "11" & x"759" => data <= x"48";
            when "11" & x"75a" => data <= x"20";
            when "11" & x"75b" => data <= x"b0";
            when "11" & x"75c" => data <= x"b4";
            when "11" & x"75d" => data <= x"68";
            when "11" & x"75e" => data <= x"90";
            when "11" & x"75f" => data <= x"95";
            when "11" & x"760" => data <= x"60";
            when "11" & x"761" => data <= x"20";
            when "11" & x"762" => data <= x"b0";
            when "11" & x"763" => data <= x"b4";
            when "11" & x"764" => data <= x"b0";
            when "11" & x"765" => data <= x"8f";
            when "11" & x"766" => data <= x"4c";
            when "11" & x"767" => data <= x"ba";
            when "11" & x"768" => data <= x"b7";
            when "11" & x"769" => data <= x"20";
            when "11" & x"76a" => data <= x"00";
            when "11" & x"76b" => data <= x"a0";
            when "11" & x"76c" => data <= x"cd";
            when "11" & x"76d" => data <= x"42";
            when "11" & x"76e" => data <= x"61";
            when "11" & x"76f" => data <= x"64";
            when "11" & x"770" => data <= x"20";
            when "11" & x"771" => data <= x"64";
            when "11" & x"772" => data <= x"72";
            when "11" & x"773" => data <= x"69";
            when "11" & x"774" => data <= x"76";
            when "11" & x"775" => data <= x"65";
            when "11" & x"776" => data <= x"00";
            when "11" & x"777" => data <= x"20";
            when "11" & x"778" => data <= x"00";
            when "11" & x"779" => data <= x"a0";
            when "11" & x"77a" => data <= x"d6";
            when "11" & x"77b" => data <= x"44";
            when "11" & x"77c" => data <= x"69";
            when "11" & x"77d" => data <= x"73";
            when "11" & x"77e" => data <= x"6b";
            when "11" & x"77f" => data <= x"20";
            when "11" & x"780" => data <= x"6e";
            when "11" & x"781" => data <= x"6f";
            when "11" & x"782" => data <= x"74";
            when "11" & x"783" => data <= x"20";
            when "11" & x"784" => data <= x"66";
            when "11" & x"785" => data <= x"6f";
            when "11" & x"786" => data <= x"75";
            when "11" & x"787" => data <= x"6e";
            when "11" & x"788" => data <= x"64";
            when "11" & x"789" => data <= x"00";
            when "11" & x"78a" => data <= x"20";
            when "11" & x"78b" => data <= x"b0";
            when "11" & x"78c" => data <= x"b4";
            when "11" & x"78d" => data <= x"b0";
            when "11" & x"78e" => data <= x"9e";
            when "11" & x"78f" => data <= x"a9";
            when "11" & x"790" => data <= x"ff";
            when "11" & x"791" => data <= x"20";
            when "11" & x"792" => data <= x"a2";
            when "11" & x"793" => data <= x"b7";
            when "11" & x"794" => data <= x"08";
            when "11" & x"795" => data <= x"e0";
            when "11" & x"796" => data <= x"04";
            when "11" & x"797" => data <= x"b0";
            when "11" & x"798" => data <= x"33";
            when "11" & x"799" => data <= x"28";
            when "11" & x"79a" => data <= x"60";
            when "11" & x"79b" => data <= x"20";
            when "11" & x"79c" => data <= x"b0";
            when "11" & x"79d" => data <= x"b4";
            when "11" & x"79e" => data <= x"b0";
            when "11" & x"79f" => data <= x"8d";
            when "11" & x"7a0" => data <= x"a5";
            when "11" & x"7a1" => data <= x"cf";
            when "11" & x"7a2" => data <= x"8d";
            when "11" & x"7a3" => data <= x"5b";
            when "11" & x"7a4" => data <= x"0d";
            when "11" & x"7a5" => data <= x"20";
            when "11" & x"7a6" => data <= x"c3";
            when "11" & x"7a7" => data <= x"b4";
            when "11" & x"7a8" => data <= x"b0";
            when "11" & x"7a9" => data <= x"26";
            when "11" & x"7aa" => data <= x"48";
            when "11" & x"7ab" => data <= x"20";
            when "11" & x"7ac" => data <= x"b0";
            when "11" & x"7ad" => data <= x"b4";
            when "11" & x"7ae" => data <= x"b0";
            when "11" & x"7af" => data <= x"15";
            when "11" & x"7b0" => data <= x"68";
            when "11" & x"7b1" => data <= x"d0";
            when "11" & x"7b2" => data <= x"b6";
            when "11" & x"7b3" => data <= x"e0";
            when "11" & x"7b4" => data <= x"04";
            when "11" & x"7b5" => data <= x"b0";
            when "11" & x"7b6" => data <= x"b2";
            when "11" & x"7b7" => data <= x"8e";
            when "11" & x"7b8" => data <= x"5b";
            when "11" & x"7b9" => data <= x"0d";
            when "11" & x"7ba" => data <= x"20";
            when "11" & x"7bb" => data <= x"c3";
            when "11" & x"7bc" => data <= x"b4";
            when "11" & x"7bd" => data <= x"b0";
            when "11" & x"7be" => data <= x"11";
            when "11" & x"7bf" => data <= x"48";
            when "11" & x"7c0" => data <= x"20";
            when "11" & x"7c1" => data <= x"b0";
            when "11" & x"7c2" => data <= x"b4";
            when "11" & x"7c3" => data <= x"90";
            when "11" & x"7c4" => data <= x"07";
            when "11" & x"7c5" => data <= x"68";
            when "11" & x"7c6" => data <= x"6a";
            when "11" & x"7c7" => data <= x"8a";
            when "11" & x"7c8" => data <= x"ae";
            when "11" & x"7c9" => data <= x"5b";
            when "11" & x"7ca" => data <= x"0d";
            when "11" & x"7cb" => data <= x"60";
            when "11" & x"7cc" => data <= x"68";
            when "11" & x"7cd" => data <= x"4c";
            when "11" & x"7ce" => data <= x"f5";
            when "11" & x"7cf" => data <= x"b6";
            when "11" & x"7d0" => data <= x"20";
            when "11" & x"7d1" => data <= x"3b";
            when "11" & x"7d2" => data <= x"b5";
            when "11" & x"7d3" => data <= x"20";
            when "11" & x"7d4" => data <= x"d7";
            when "11" & x"7d5" => data <= x"b1";
            when "11" & x"7d6" => data <= x"ad";
            when "11" & x"7d7" => data <= x"5c";
            when "11" & x"7d8" => data <= x"0d";
            when "11" & x"7d9" => data <= x"f0";
            when "11" & x"7da" => data <= x"f2";
            when "11" & x"7db" => data <= x"ad";
            when "11" & x"7dc" => data <= x"5e";
            when "11" & x"7dd" => data <= x"0d";
            when "11" & x"7de" => data <= x"d0";
            when "11" & x"7df" => data <= x"ed";
            when "11" & x"7e0" => data <= x"ad";
            when "11" & x"7e1" => data <= x"54";
            when "11" & x"7e2" => data <= x"0d";
            when "11" & x"7e3" => data <= x"30";
            when "11" & x"7e4" => data <= x"92";
            when "11" & x"7e5" => data <= x"20";
            when "11" & x"7e6" => data <= x"b3";
            when "11" & x"7e7" => data <= x"b5";
            when "11" & x"7e8" => data <= x"90";
            when "11" & x"7e9" => data <= x"06";
            when "11" & x"7ea" => data <= x"20";
            when "11" & x"7eb" => data <= x"fc";
            when "11" & x"7ec" => data <= x"b1";
            when "11" & x"7ed" => data <= x"4c";
            when "11" & x"7ee" => data <= x"e0";
            when "11" & x"7ef" => data <= x"b7";
            when "11" & x"7f0" => data <= x"ad";
            when "11" & x"7f1" => data <= x"54";
            when "11" & x"7f2" => data <= x"0d";
            when "11" & x"7f3" => data <= x"6a";
            when "11" & x"7f4" => data <= x"ad";
            when "11" & x"7f5" => data <= x"53";
            when "11" & x"7f6" => data <= x"0d";
            when "11" & x"7f7" => data <= x"ae";
            when "11" & x"7f8" => data <= x"5b";
            when "11" & x"7f9" => data <= x"0d";
            when "11" & x"7fa" => data <= x"60";
            when "11" & x"7fb" => data <= x"20";
            when "11" & x"7fc" => data <= x"61";
            when "11" & x"7fd" => data <= x"b7";
            when "11" & x"7fe" => data <= x"a6";
            when "11" & x"7ff" => data <= x"cf";
            when "11" & x"800" => data <= x"20";
            when "11" & x"801" => data <= x"0f";
            when "11" & x"802" => data <= x"b0";
            when "11" & x"803" => data <= x"4c";
            when "11" & x"804" => data <= x"07";
            when "11" & x"805" => data <= x"94";
            when "11" & x"806" => data <= x"20";
            when "11" & x"807" => data <= x"9b";
            when "11" & x"808" => data <= x"b7";
            when "11" & x"809" => data <= x"4c";
            when "11" & x"80a" => data <= x"0f";
            when "11" & x"80b" => data <= x"b0";
            when "11" & x"80c" => data <= x"a9";
            when "11" & x"80d" => data <= x"00";
            when "11" & x"80e" => data <= x"8d";
            when "11" & x"80f" => data <= x"57";
            when "11" & x"810" => data <= x"0d";
            when "11" & x"811" => data <= x"8d";
            when "11" & x"812" => data <= x"58";
            when "11" & x"813" => data <= x"0d";
            when "11" & x"814" => data <= x"20";
            when "11" & x"815" => data <= x"c3";
            when "11" & x"816" => data <= x"b4";
            when "11" & x"817" => data <= x"b0";
            when "11" & x"818" => data <= x"2d";
            when "11" & x"819" => data <= x"8e";
            when "11" & x"81a" => data <= x"59";
            when "11" & x"81b" => data <= x"0d";
            when "11" & x"81c" => data <= x"8e";
            when "11" & x"81d" => data <= x"53";
            when "11" & x"81e" => data <= x"0d";
            when "11" & x"81f" => data <= x"8d";
            when "11" & x"820" => data <= x"5a";
            when "11" & x"821" => data <= x"0d";
            when "11" & x"822" => data <= x"8d";
            when "11" & x"823" => data <= x"54";
            when "11" & x"824" => data <= x"0d";
            when "11" & x"825" => data <= x"20";
            when "11" & x"826" => data <= x"c3";
            when "11" & x"827" => data <= x"b4";
            when "11" & x"828" => data <= x"b0";
            when "11" & x"829" => data <= x"25";
            when "11" & x"82a" => data <= x"8e";
            when "11" & x"82b" => data <= x"59";
            when "11" & x"82c" => data <= x"0d";
            when "11" & x"82d" => data <= x"8d";
            when "11" & x"82e" => data <= x"5a";
            when "11" & x"82f" => data <= x"0d";
            when "11" & x"830" => data <= x"ec";
            when "11" & x"831" => data <= x"53";
            when "11" & x"832" => data <= x"0d";
            when "11" & x"833" => data <= x"ed";
            when "11" & x"834" => data <= x"54";
            when "11" & x"835" => data <= x"0d";
            when "11" & x"836" => data <= x"10";
            when "11" & x"837" => data <= x"1f";
            when "11" & x"838" => data <= x"20";
            when "11" & x"839" => data <= x"00";
            when "11" & x"83a" => data <= x"a0";
            when "11" & x"83b" => data <= x"ff";
            when "11" & x"83c" => data <= x"42";
            when "11" & x"83d" => data <= x"61";
            when "11" & x"83e" => data <= x"64";
            when "11" & x"83f" => data <= x"20";
            when "11" & x"840" => data <= x"72";
            when "11" & x"841" => data <= x"61";
            when "11" & x"842" => data <= x"6e";
            when "11" & x"843" => data <= x"67";
            when "11" & x"844" => data <= x"65";
            when "11" & x"845" => data <= x"00";
            when "11" & x"846" => data <= x"a2";
            when "11" & x"847" => data <= x"fe";
            when "11" & x"848" => data <= x"8e";
            when "11" & x"849" => data <= x"59";
            when "11" & x"84a" => data <= x"0d";
            when "11" & x"84b" => data <= x"e8";
            when "11" & x"84c" => data <= x"8e";
            when "11" & x"84d" => data <= x"5a";
            when "11" & x"84e" => data <= x"0d";
            when "11" & x"84f" => data <= x"a9";
            when "11" & x"850" => data <= x"00";
            when "11" & x"851" => data <= x"8d";
            when "11" & x"852" => data <= x"53";
            when "11" & x"853" => data <= x"0d";
            when "11" & x"854" => data <= x"8d";
            when "11" & x"855" => data <= x"54";
            when "11" & x"856" => data <= x"0d";
            when "11" & x"857" => data <= x"ee";
            when "11" & x"858" => data <= x"59";
            when "11" & x"859" => data <= x"0d";
            when "11" & x"85a" => data <= x"d0";
            when "11" & x"85b" => data <= x"03";
            when "11" & x"85c" => data <= x"ee";
            when "11" & x"85d" => data <= x"5a";
            when "11" & x"85e" => data <= x"0d";
            when "11" & x"85f" => data <= x"20";
            when "11" & x"860" => data <= x"3b";
            when "11" & x"861" => data <= x"b5";
            when "11" & x"862" => data <= x"ad";
            when "11" & x"863" => data <= x"54";
            when "11" & x"864" => data <= x"0d";
            when "11" & x"865" => data <= x"6a";
            when "11" & x"866" => data <= x"ad";
            when "11" & x"867" => data <= x"53";
            when "11" & x"868" => data <= x"0d";
            when "11" & x"869" => data <= x"20";
            when "11" & x"86a" => data <= x"a0";
            when "11" & x"86b" => data <= x"b1";
            when "11" & x"86c" => data <= x"a2";
            when "11" & x"86d" => data <= x"00";
            when "11" & x"86e" => data <= x"ad";
            when "11" & x"86f" => data <= x"5c";
            when "11" & x"870" => data <= x"0d";
            when "11" & x"871" => data <= x"d0";
            when "11" & x"872" => data <= x"04";
            when "11" & x"873" => data <= x"ca";
            when "11" & x"874" => data <= x"8e";
            when "11" & x"875" => data <= x"5e";
            when "11" & x"876" => data <= x"0d";
            when "11" & x"877" => data <= x"ad";
            when "11" & x"878" => data <= x"54";
            when "11" & x"879" => data <= x"0d";
            when "11" & x"87a" => data <= x"30";
            when "11" & x"87b" => data <= x"33";
            when "11" & x"87c" => data <= x"ad";
            when "11" & x"87d" => data <= x"53";
            when "11" & x"87e" => data <= x"0d";
            when "11" & x"87f" => data <= x"cd";
            when "11" & x"880" => data <= x"59";
            when "11" & x"881" => data <= x"0d";
            when "11" & x"882" => data <= x"ad";
            when "11" & x"883" => data <= x"54";
            when "11" & x"884" => data <= x"0d";
            when "11" & x"885" => data <= x"ed";
            when "11" & x"886" => data <= x"5a";
            when "11" & x"887" => data <= x"0d";
            when "11" & x"888" => data <= x"b0";
            when "11" & x"889" => data <= x"25";
            when "11" & x"88a" => data <= x"20";
            when "11" & x"88b" => data <= x"b3";
            when "11" & x"88c" => data <= x"b5";
            when "11" & x"88d" => data <= x"b0";
            when "11" & x"88e" => data <= x"16";
            when "11" & x"88f" => data <= x"20";
            when "11" & x"890" => data <= x"e5";
            when "11" & x"891" => data <= x"b5";
            when "11" & x"892" => data <= x"f8";
            when "11" & x"893" => data <= x"18";
            when "11" & x"894" => data <= x"ad";
            when "11" & x"895" => data <= x"57";
            when "11" & x"896" => data <= x"0d";
            when "11" & x"897" => data <= x"69";
            when "11" & x"898" => data <= x"01";
            when "11" & x"899" => data <= x"8d";
            when "11" & x"89a" => data <= x"57";
            when "11" & x"89b" => data <= x"0d";
            when "11" & x"89c" => data <= x"ad";
            when "11" & x"89d" => data <= x"58";
            when "11" & x"89e" => data <= x"0d";
            when "11" & x"89f" => data <= x"69";
            when "11" & x"8a0" => data <= x"00";
            when "11" & x"8a1" => data <= x"8d";
            when "11" & x"8a2" => data <= x"58";
            when "11" & x"8a3" => data <= x"0d";
            when "11" & x"8a4" => data <= x"d8";
            when "11" & x"8a5" => data <= x"24";
            when "11" & x"8a6" => data <= x"ff";
            when "11" & x"8a7" => data <= x"30";
            when "11" & x"8a8" => data <= x"47";
            when "11" & x"8a9" => data <= x"20";
            when "11" & x"8aa" => data <= x"fc";
            when "11" & x"8ab" => data <= x"b1";
            when "11" & x"8ac" => data <= x"4c";
            when "11" & x"8ad" => data <= x"77";
            when "11" & x"8ae" => data <= x"b8";
            when "11" & x"8af" => data <= x"a9";
            when "11" & x"8b0" => data <= x"86";
            when "11" & x"8b1" => data <= x"20";
            when "11" & x"8b2" => data <= x"f4";
            when "11" & x"8b3" => data <= x"ff";
            when "11" & x"8b4" => data <= x"e0";
            when "11" & x"8b5" => data <= x"00";
            when "11" & x"8b6" => data <= x"f0";
            when "11" & x"8b7" => data <= x"03";
            when "11" & x"8b8" => data <= x"20";
            when "11" & x"8b9" => data <= x"e7";
            when "11" & x"8ba" => data <= x"ff";
            when "11" & x"8bb" => data <= x"ad";
            when "11" & x"8bc" => data <= x"58";
            when "11" & x"8bd" => data <= x"0d";
            when "11" & x"8be" => data <= x"a2";
            when "11" & x"8bf" => data <= x"00";
            when "11" & x"8c0" => data <= x"a0";
            when "11" & x"8c1" => data <= x"04";
            when "11" & x"8c2" => data <= x"20";
            when "11" & x"8c3" => data <= x"26";
            when "11" & x"8c4" => data <= x"b6";
            when "11" & x"8c5" => data <= x"ad";
            when "11" & x"8c6" => data <= x"57";
            when "11" & x"8c7" => data <= x"0d";
            when "11" & x"8c8" => data <= x"20";
            when "11" & x"8c9" => data <= x"26";
            when "11" & x"8ca" => data <= x"b6";
            when "11" & x"8cb" => data <= x"20";
            when "11" & x"8cc" => data <= x"44";
            when "11" & x"8cd" => data <= x"b6";
            when "11" & x"8ce" => data <= x"20";
            when "11" & x"8cf" => data <= x"64";
            when "11" & x"8d0" => data <= x"69";
            when "11" & x"8d1" => data <= x"73";
            when "11" & x"8d2" => data <= x"6b";
            when "11" & x"8d3" => data <= x"00";
            when "11" & x"8d4" => data <= x"ad";
            when "11" & x"8d5" => data <= x"58";
            when "11" & x"8d6" => data <= x"0d";
            when "11" & x"8d7" => data <= x"d0";
            when "11" & x"8d8" => data <= x"05";
            when "11" & x"8d9" => data <= x"ce";
            when "11" & x"8da" => data <= x"57";
            when "11" & x"8db" => data <= x"0d";
            when "11" & x"8dc" => data <= x"f0";
            when "11" & x"8dd" => data <= x"05";
            when "11" & x"8de" => data <= x"a9";
            when "11" & x"8df" => data <= x"73";
            when "11" & x"8e0" => data <= x"20";
            when "11" & x"8e1" => data <= x"ee";
            when "11" & x"8e2" => data <= x"ff";
            when "11" & x"8e3" => data <= x"20";
            when "11" & x"8e4" => data <= x"44";
            when "11" & x"8e5" => data <= x"b6";
            when "11" & x"8e6" => data <= x"20";
            when "11" & x"8e7" => data <= x"66";
            when "11" & x"8e8" => data <= x"6f";
            when "11" & x"8e9" => data <= x"75";
            when "11" & x"8ea" => data <= x"6e";
            when "11" & x"8eb" => data <= x"64";
            when "11" & x"8ec" => data <= x"00";
            when "11" & x"8ed" => data <= x"4c";
            when "11" & x"8ee" => data <= x"e7";
            when "11" & x"8ef" => data <= x"ff";
            when "11" & x"8f0" => data <= x"4c";
            when "11" & x"8f1" => data <= x"82";
            when "11" & x"8f2" => data <= x"a0";
            when "11" & x"8f3" => data <= x"4c";
            when "11" & x"8f4" => data <= x"f5";
            when "11" & x"8f5" => data <= x"b6";
            when "11" & x"8f6" => data <= x"20";
            when "11" & x"8f7" => data <= x"b0";
            when "11" & x"8f8" => data <= x"b4";
            when "11" & x"8f9" => data <= x"90";
            when "11" & x"8fa" => data <= x"f8";
            when "11" & x"8fb" => data <= x"a2";
            when "11" & x"8fc" => data <= x"00";
            when "11" & x"8fd" => data <= x"8e";
            when "11" & x"8fe" => data <= x"57";
            when "11" & x"8ff" => data <= x"0d";
            when "11" & x"900" => data <= x"8e";
            when "11" & x"901" => data <= x"58";
            when "11" & x"902" => data <= x"0d";
            when "11" & x"903" => data <= x"8e";
            when "11" & x"904" => data <= x"59";
            when "11" & x"905" => data <= x"0d";
            when "11" & x"906" => data <= x"8e";
            when "11" & x"907" => data <= x"5a";
            when "11" & x"908" => data <= x"0d";
            when "11" & x"909" => data <= x"a9";
            when "11" & x"90a" => data <= x"80";
            when "11" & x"90b" => data <= x"20";
            when "11" & x"90c" => data <= x"9c";
            when "11" & x"90d" => data <= x"b0";
            when "11" & x"90e" => data <= x"a9";
            when "11" & x"90f" => data <= x"10";
            when "11" & x"910" => data <= x"85";
            when "11" & x"911" => data <= x"f2";
            when "11" & x"912" => data <= x"a9";
            when "11" & x"913" => data <= x"0e";
            when "11" & x"914" => data <= x"85";
            when "11" & x"915" => data <= x"f3";
            when "11" & x"916" => data <= x"a0";
            when "11" & x"917" => data <= x"0f";
            when "11" & x"918" => data <= x"b1";
            when "11" & x"919" => data <= x"f2";
            when "11" & x"91a" => data <= x"c9";
            when "11" & x"91b" => data <= x"ff";
            when "11" & x"91c" => data <= x"f0";
            when "11" & x"91d" => data <= x"42";
            when "11" & x"91e" => data <= x"f8";
            when "11" & x"91f" => data <= x"a8";
            when "11" & x"920" => data <= x"10";
            when "11" & x"921" => data <= x"0e";
            when "11" & x"922" => data <= x"18";
            when "11" & x"923" => data <= x"ad";
            when "11" & x"924" => data <= x"57";
            when "11" & x"925" => data <= x"0d";
            when "11" & x"926" => data <= x"69";
            when "11" & x"927" => data <= x"01";
            when "11" & x"928" => data <= x"8d";
            when "11" & x"929" => data <= x"57";
            when "11" & x"92a" => data <= x"0d";
            when "11" & x"92b" => data <= x"90";
            when "11" & x"92c" => data <= x"03";
            when "11" & x"92d" => data <= x"ee";
            when "11" & x"92e" => data <= x"58";
            when "11" & x"92f" => data <= x"0d";
            when "11" & x"930" => data <= x"18";
            when "11" & x"931" => data <= x"ad";
            when "11" & x"932" => data <= x"59";
            when "11" & x"933" => data <= x"0d";
            when "11" & x"934" => data <= x"69";
            when "11" & x"935" => data <= x"01";
            when "11" & x"936" => data <= x"8d";
            when "11" & x"937" => data <= x"59";
            when "11" & x"938" => data <= x"0d";
            when "11" & x"939" => data <= x"90";
            when "11" & x"93a" => data <= x"03";
            when "11" & x"93b" => data <= x"ee";
            when "11" & x"93c" => data <= x"5a";
            when "11" & x"93d" => data <= x"0d";
            when "11" & x"93e" => data <= x"d8";
            when "11" & x"93f" => data <= x"18";
            when "11" & x"940" => data <= x"a5";
            when "11" & x"941" => data <= x"f2";
            when "11" & x"942" => data <= x"69";
            when "11" & x"943" => data <= x"10";
            when "11" & x"944" => data <= x"85";
            when "11" & x"945" => data <= x"f2";
            when "11" & x"946" => data <= x"d0";
            when "11" & x"947" => data <= x"ce";
            when "11" & x"948" => data <= x"a5";
            when "11" & x"949" => data <= x"f3";
            when "11" & x"94a" => data <= x"49";
            when "11" & x"94b" => data <= x"01";
            when "11" & x"94c" => data <= x"85";
            when "11" & x"94d" => data <= x"f3";
            when "11" & x"94e" => data <= x"6a";
            when "11" & x"94f" => data <= x"b0";
            when "11" & x"950" => data <= x"c5";
            when "11" & x"951" => data <= x"ad";
            when "11" & x"952" => data <= x"82";
            when "11" & x"953" => data <= x"10";
            when "11" & x"954" => data <= x"69";
            when "11" & x"955" => data <= x"01";
            when "11" & x"956" => data <= x"c9";
            when "11" & x"957" => data <= x"90";
            when "11" & x"958" => data <= x"f0";
            when "11" & x"959" => data <= x"06";
            when "11" & x"95a" => data <= x"20";
            when "11" & x"95b" => data <= x"9c";
            when "11" & x"95c" => data <= x"b0";
            when "11" & x"95d" => data <= x"4c";
            when "11" & x"95e" => data <= x"16";
            when "11" & x"95f" => data <= x"b9";
            when "11" & x"960" => data <= x"a0";
            when "11" & x"961" => data <= x"04";
            when "11" & x"962" => data <= x"a2";
            when "11" & x"963" => data <= x"00";
            when "11" & x"964" => data <= x"ad";
            when "11" & x"965" => data <= x"58";
            when "11" & x"966" => data <= x"0d";
            when "11" & x"967" => data <= x"20";
            when "11" & x"968" => data <= x"26";
            when "11" & x"969" => data <= x"b6";
            when "11" & x"96a" => data <= x"ad";
            when "11" & x"96b" => data <= x"57";
            when "11" & x"96c" => data <= x"0d";
            when "11" & x"96d" => data <= x"20";
            when "11" & x"96e" => data <= x"26";
            when "11" & x"96f" => data <= x"b6";
            when "11" & x"970" => data <= x"20";
            when "11" & x"971" => data <= x"44";
            when "11" & x"972" => data <= x"b6";
            when "11" & x"973" => data <= x"20";
            when "11" & x"974" => data <= x"6f";
            when "11" & x"975" => data <= x"66";
            when "11" & x"976" => data <= x"20";
            when "11" & x"977" => data <= x"00";
            when "11" & x"978" => data <= x"a2";
            when "11" & x"979" => data <= x"00";
            when "11" & x"97a" => data <= x"a0";
            when "11" & x"97b" => data <= x"04";
            when "11" & x"97c" => data <= x"ad";
            when "11" & x"97d" => data <= x"5a";
            when "11" & x"97e" => data <= x"0d";
            when "11" & x"97f" => data <= x"20";
            when "11" & x"980" => data <= x"26";
            when "11" & x"981" => data <= x"b6";
            when "11" & x"982" => data <= x"ad";
            when "11" & x"983" => data <= x"59";
            when "11" & x"984" => data <= x"0d";
            when "11" & x"985" => data <= x"20";
            when "11" & x"986" => data <= x"26";
            when "11" & x"987" => data <= x"b6";
            when "11" & x"988" => data <= x"20";
            when "11" & x"989" => data <= x"44";
            when "11" & x"98a" => data <= x"b6";
            when "11" & x"98b" => data <= x"20";
            when "11" & x"98c" => data <= x"64";
            when "11" & x"98d" => data <= x"69";
            when "11" & x"98e" => data <= x"73";
            when "11" & x"98f" => data <= x"6b";
            when "11" & x"990" => data <= x"00";
            when "11" & x"991" => data <= x"ad";
            when "11" & x"992" => data <= x"5a";
            when "11" & x"993" => data <= x"0d";
            when "11" & x"994" => data <= x"d0";
            when "11" & x"995" => data <= x"07";
            when "11" & x"996" => data <= x"ad";
            when "11" & x"997" => data <= x"59";
            when "11" & x"998" => data <= x"0d";
            when "11" & x"999" => data <= x"c9";
            when "11" & x"99a" => data <= x"01";
            when "11" & x"99b" => data <= x"f0";
            when "11" & x"99c" => data <= x"05";
            when "11" & x"99d" => data <= x"a9";
            when "11" & x"99e" => data <= x"73";
            when "11" & x"99f" => data <= x"20";
            when "11" & x"9a0" => data <= x"ee";
            when "11" & x"9a1" => data <= x"ff";
            when "11" & x"9a2" => data <= x"20";
            when "11" & x"9a3" => data <= x"44";
            when "11" & x"9a4" => data <= x"b6";
            when "11" & x"9a5" => data <= x"20";
            when "11" & x"9a6" => data <= x"66";
            when "11" & x"9a7" => data <= x"72";
            when "11" & x"9a8" => data <= x"65";
            when "11" & x"9a9" => data <= x"65";
            when "11" & x"9aa" => data <= x"20";
            when "11" & x"9ab" => data <= x"28";
            when "11" & x"9ac" => data <= x"75";
            when "11" & x"9ad" => data <= x"6e";
            when "11" & x"9ae" => data <= x"66";
            when "11" & x"9af" => data <= x"6f";
            when "11" & x"9b0" => data <= x"72";
            when "11" & x"9b1" => data <= x"6d";
            when "11" & x"9b2" => data <= x"61";
            when "11" & x"9b3" => data <= x"74";
            when "11" & x"9b4" => data <= x"74";
            when "11" & x"9b5" => data <= x"65";
            when "11" & x"9b6" => data <= x"64";
            when "11" & x"9b7" => data <= x"29";
            when "11" & x"9b8" => data <= x"00";
            when "11" & x"9b9" => data <= x"4c";
            when "11" & x"9ba" => data <= x"e7";
            when "11" & x"9bb" => data <= x"ff";
            when "11" & x"9bc" => data <= x"20";
            when "11" & x"9bd" => data <= x"30";
            when "11" & x"9be" => data <= x"b7";
            when "11" & x"9bf" => data <= x"a2";
            when "11" & x"9c0" => data <= x"04";
            when "11" & x"9c1" => data <= x"8e";
            when "11" & x"9c2" => data <= x"5b";
            when "11" & x"9c3" => data <= x"0d";
            when "11" & x"9c4" => data <= x"a2";
            when "11" & x"9c5" => data <= x"00";
            when "11" & x"9c6" => data <= x"b0";
            when "11" & x"9c7" => data <= x"06";
            when "11" & x"9c8" => data <= x"aa";
            when "11" & x"9c9" => data <= x"e8";
            when "11" & x"9ca" => data <= x"8e";
            when "11" & x"9cb" => data <= x"5b";
            when "11" & x"9cc" => data <= x"0d";
            when "11" & x"9cd" => data <= x"ca";
            when "11" & x"9ce" => data <= x"8a";
            when "11" & x"9cf" => data <= x"48";
            when "11" & x"9d0" => data <= x"a2";
            when "11" & x"9d1" => data <= x"20";
            when "11" & x"9d2" => data <= x"a0";
            when "11" & x"9d3" => data <= x"02";
            when "11" & x"9d4" => data <= x"20";
            when "11" & x"9d5" => data <= x"26";
            when "11" & x"9d6" => data <= x"b6";
            when "11" & x"9d7" => data <= x"a9";
            when "11" & x"9d8" => data <= x"3a";
            when "11" & x"9d9" => data <= x"20";
            when "11" & x"9da" => data <= x"ee";
            when "11" & x"9db" => data <= x"ff";
            when "11" & x"9dc" => data <= x"68";
            when "11" & x"9dd" => data <= x"aa";
            when "11" & x"9de" => data <= x"48";
            when "11" & x"9df" => data <= x"bd";
            when "11" & x"9e0" => data <= x"10";
            when "11" & x"9e1" => data <= x"0d";
            when "11" & x"9e2" => data <= x"30";
            when "11" & x"9e3" => data <= x"0f";
            when "11" & x"9e4" => data <= x"6a";
            when "11" & x"9e5" => data <= x"bd";
            when "11" & x"9e6" => data <= x"0c";
            when "11" & x"9e7" => data <= x"0d";
            when "11" & x"9e8" => data <= x"20";
            when "11" & x"9e9" => data <= x"a0";
            when "11" & x"9ea" => data <= x"b1";
            when "11" & x"9eb" => data <= x"c9";
            when "11" & x"9ec" => data <= x"ff";
            when "11" & x"9ed" => data <= x"f0";
            when "11" & x"9ee" => data <= x"04";
            when "11" & x"9ef" => data <= x"38";
            when "11" & x"9f0" => data <= x"20";
            when "11" & x"9f1" => data <= x"e5";
            when "11" & x"9f2" => data <= x"b5";
            when "11" & x"9f3" => data <= x"20";
            when "11" & x"9f4" => data <= x"e7";
            when "11" & x"9f5" => data <= x"ff";
            when "11" & x"9f6" => data <= x"68";
            when "11" & x"9f7" => data <= x"aa";
            when "11" & x"9f8" => data <= x"e8";
            when "11" & x"9f9" => data <= x"ec";
            when "11" & x"9fa" => data <= x"5b";
            when "11" & x"9fb" => data <= x"0d";
            when "11" & x"9fc" => data <= x"90";
            when "11" & x"9fd" => data <= x"d0";
            when "11" & x"9fe" => data <= x"60";
            when "11" & x"9ff" => data <= x"4c";
            when "11" & x"a00" => data <= x"f5";
            when "11" & x"a01" => data <= x"b6";
            when "11" & x"a02" => data <= x"a9";
            when "11" & x"a03" => data <= x"00";
            when "11" & x"a04" => data <= x"f0";
            when "11" & x"a05" => data <= x"02";
            when "11" & x"a06" => data <= x"a9";
            when "11" & x"a07" => data <= x"0f";
            when "11" & x"a08" => data <= x"48";
            when "11" & x"a09" => data <= x"20";
            when "11" & x"a0a" => data <= x"61";
            when "11" & x"a0b" => data <= x"b7";
            when "11" & x"a0c" => data <= x"20";
            when "11" & x"a0d" => data <= x"c1";
            when "11" & x"a0e" => data <= x"af";
            when "11" & x"a0f" => data <= x"30";
            when "11" & x"a10" => data <= x"0e";
            when "11" & x"a11" => data <= x"68";
            when "11" & x"a12" => data <= x"b0";
            when "11" & x"a13" => data <= x"05";
            when "11" & x"a14" => data <= x"99";
            when "11" & x"a15" => data <= x"00";
            when "11" & x"a16" => data <= x"0e";
            when "11" & x"a17" => data <= x"90";
            when "11" & x"a18" => data <= x"03";
            when "11" & x"a19" => data <= x"99";
            when "11" & x"a1a" => data <= x"00";
            when "11" & x"a1b" => data <= x"0f";
            when "11" & x"a1c" => data <= x"4c";
            when "11" & x"a1d" => data <= x"cd";
            when "11" & x"a1e" => data <= x"b0";
            when "11" & x"a1f" => data <= x"c9";
            when "11" & x"a20" => data <= x"ff";
            when "11" & x"a21" => data <= x"f0";
            when "11" & x"a22" => data <= x"03";
            when "11" & x"a23" => data <= x"4c";
            when "11" & x"a24" => data <= x"59";
            when "11" & x"a25" => data <= x"b0";
            when "11" & x"a26" => data <= x"4c";
            when "11" & x"a27" => data <= x"3f";
            when "11" & x"a28" => data <= x"b0";
            when "11" & x"a29" => data <= x"20";
            when "11" & x"a2a" => data <= x"bd";
            when "11" & x"a2b" => data <= x"9b";
            when "11" & x"a2c" => data <= x"20";
            when "11" & x"a2d" => data <= x"4f";
            when "11" & x"a2e" => data <= x"b7";
            when "11" & x"a2f" => data <= x"6a";
            when "11" & x"a30" => data <= x"08";
            when "11" & x"a31" => data <= x"8a";
            when "11" & x"a32" => data <= x"48";
            when "11" & x"a33" => data <= x"20";
            when "11" & x"a34" => data <= x"c1";
            when "11" & x"a35" => data <= x"af";
            when "11" & x"a36" => data <= x"30";
            when "11" & x"a37" => data <= x"e7";
            when "11" & x"a38" => data <= x"68";
            when "11" & x"a39" => data <= x"28";
            when "11" & x"a3a" => data <= x"20";
            when "11" & x"a3b" => data <= x"a0";
            when "11" & x"a3c" => data <= x"b1";
            when "11" & x"a3d" => data <= x"20";
            when "11" & x"a3e" => data <= x"44";
            when "11" & x"a3f" => data <= x"b6";
            when "11" & x"a40" => data <= x"4b";
            when "11" & x"a41" => data <= x"69";
            when "11" & x"a42" => data <= x"6c";
            when "11" & x"a43" => data <= x"6c";
            when "11" & x"a44" => data <= x"00";
            when "11" & x"a45" => data <= x"38";
            when "11" & x"a46" => data <= x"20";
            when "11" & x"a47" => data <= x"e5";
            when "11" & x"a48" => data <= x"b5";
            when "11" & x"a49" => data <= x"20";
            when "11" & x"a4a" => data <= x"44";
            when "11" & x"a4b" => data <= x"b6";
            when "11" & x"a4c" => data <= x"20";
            when "11" & x"a4d" => data <= x"3a";
            when "11" & x"a4e" => data <= x"20";
            when "11" & x"a4f" => data <= x"00";
            when "11" & x"a50" => data <= x"20";
            when "11" & x"a51" => data <= x"9e";
            when "11" & x"a52" => data <= x"9c";
            when "11" & x"a53" => data <= x"08";
            when "11" & x"a54" => data <= x"20";
            when "11" & x"a55" => data <= x"e7";
            when "11" & x"a56" => data <= x"ff";
            when "11" & x"a57" => data <= x"28";
            when "11" & x"a58" => data <= x"d0";
            when "11" & x"a59" => data <= x"09";
            when "11" & x"a5a" => data <= x"a0";
            when "11" & x"a5b" => data <= x"0f";
            when "11" & x"a5c" => data <= x"a9";
            when "11" & x"a5d" => data <= x"f0";
            when "11" & x"a5e" => data <= x"91";
            when "11" & x"a5f" => data <= x"f2";
            when "11" & x"a60" => data <= x"4c";
            when "11" & x"a61" => data <= x"cd";
            when "11" & x"a62" => data <= x"b0";
            when "11" & x"a63" => data <= x"60";
            when "11" & x"a64" => data <= x"a9";
            when "11" & x"a65" => data <= x"00";
            when "11" & x"a66" => data <= x"20";
            when "11" & x"a67" => data <= x"6e";
            when "11" & x"a68" => data <= x"ba";
            when "11" & x"a69" => data <= x"4c";
            when "11" & x"a6a" => data <= x"63";
            when "11" & x"a6b" => data <= x"af";
            when "11" & x"a6c" => data <= x"a9";
            when "11" & x"a6d" => data <= x"01";
            when "11" & x"a6e" => data <= x"8d";
            when "11" & x"a6f" => data <= x"5f";
            when "11" & x"a70" => data <= x"0d";
            when "11" & x"a71" => data <= x"20";
            when "11" & x"a72" => data <= x"4f";
            when "11" & x"a73" => data <= x"b7";
            when "11" & x"a74" => data <= x"6a";
            when "11" & x"a75" => data <= x"08";
            when "11" & x"a76" => data <= x"8a";
            when "11" & x"a77" => data <= x"48";
            when "11" & x"a78" => data <= x"20";
            when "11" & x"a79" => data <= x"c1";
            when "11" & x"a7a" => data <= x"af";
            when "11" & x"a7b" => data <= x"10";
            when "11" & x"a7c" => data <= x"26";
            when "11" & x"a7d" => data <= x"aa";
            when "11" & x"a7e" => data <= x"e8";
            when "11" & x"a7f" => data <= x"f0";
            when "11" & x"a80" => data <= x"3d";
            when "11" & x"a81" => data <= x"98";
            when "11" & x"a82" => data <= x"29";
            when "11" & x"a83" => data <= x"f0";
            when "11" & x"a84" => data <= x"85";
            when "11" & x"a85" => data <= x"f2";
            when "11" & x"a86" => data <= x"a0";
            when "11" & x"a87" => data <= x"0e";
            when "11" & x"a88" => data <= x"90";
            when "11" & x"a89" => data <= x"01";
            when "11" & x"a8a" => data <= x"c8";
            when "11" & x"a8b" => data <= x"84";
            when "11" & x"a8c" => data <= x"f3";
            when "11" & x"a8d" => data <= x"a0";
            when "11" & x"a8e" => data <= x"0f";
            when "11" & x"a8f" => data <= x"98";
            when "11" & x"a90" => data <= x"91";
            when "11" & x"a91" => data <= x"f2";
            when "11" & x"a92" => data <= x"ad";
            when "11" & x"a93" => data <= x"5f";
            when "11" & x"a94" => data <= x"0d";
            when "11" & x"a95" => data <= x"d0";
            when "11" & x"a96" => data <= x"06";
            when "11" & x"a97" => data <= x"88";
            when "11" & x"a98" => data <= x"91";
            when "11" & x"a99" => data <= x"f2";
            when "11" & x"a9a" => data <= x"88";
            when "11" & x"a9b" => data <= x"10";
            when "11" & x"a9c" => data <= x"fb";
            when "11" & x"a9d" => data <= x"20";
            when "11" & x"a9e" => data <= x"cd";
            when "11" & x"a9f" => data <= x"b0";
            when "11" & x"aa0" => data <= x"68";
            when "11" & x"aa1" => data <= x"28";
            when "11" & x"aa2" => data <= x"60";
            when "11" & x"aa3" => data <= x"20";
            when "11" & x"aa4" => data <= x"00";
            when "11" & x"aa5" => data <= x"a0";
            when "11" & x"aa6" => data <= x"ff";
            when "11" & x"aa7" => data <= x"44";
            when "11" & x"aa8" => data <= x"69";
            when "11" & x"aa9" => data <= x"73";
            when "11" & x"aaa" => data <= x"6b";
            when "11" & x"aab" => data <= x"20";
            when "11" & x"aac" => data <= x"61";
            when "11" & x"aad" => data <= x"6c";
            when "11" & x"aae" => data <= x"72";
            when "11" & x"aaf" => data <= x"65";
            when "11" & x"ab0" => data <= x"61";
            when "11" & x"ab1" => data <= x"64";
            when "11" & x"ab2" => data <= x"79";
            when "11" & x"ab3" => data <= x"20";
            when "11" & x"ab4" => data <= x"66";
            when "11" & x"ab5" => data <= x"6f";
            when "11" & x"ab6" => data <= x"72";
            when "11" & x"ab7" => data <= x"6d";
            when "11" & x"ab8" => data <= x"61";
            when "11" & x"ab9" => data <= x"74";
            when "11" & x"aba" => data <= x"74";
            when "11" & x"abb" => data <= x"65";
            when "11" & x"abc" => data <= x"64";
            when "11" & x"abd" => data <= x"00";
            when "11" & x"abe" => data <= x"4c";
            when "11" & x"abf" => data <= x"3f";
            when "11" & x"ac0" => data <= x"b0";
            when "11" & x"ac1" => data <= x"20";
            when "11" & x"ac2" => data <= x"30";
            when "11" & x"ac3" => data <= x"b7";
            when "11" & x"ac4" => data <= x"8d";
            when "11" & x"ac5" => data <= x"5b";
            when "11" & x"ac6" => data <= x"0d";
            when "11" & x"ac7" => data <= x"20";
            when "11" & x"ac8" => data <= x"25";
            when "11" & x"ac9" => data <= x"bb";
            when "11" & x"aca" => data <= x"08";
            when "11" & x"acb" => data <= x"48";
            when "11" & x"acc" => data <= x"a9";
            when "11" & x"acd" => data <= x"0f";
            when "11" & x"ace" => data <= x"91";
            when "11" & x"acf" => data <= x"f2";
            when "11" & x"ad0" => data <= x"88";
            when "11" & x"ad1" => data <= x"a9";
            when "11" & x"ad2" => data <= x"00";
            when "11" & x"ad3" => data <= x"91";
            when "11" & x"ad4" => data <= x"f2";
            when "11" & x"ad5" => data <= x"88";
            when "11" & x"ad6" => data <= x"10";
            when "11" & x"ad7" => data <= x"fb";
            when "11" & x"ad8" => data <= x"20";
            when "11" & x"ad9" => data <= x"b8";
            when "11" & x"ada" => data <= x"b0";
            when "11" & x"adb" => data <= x"68";
            when "11" & x"adc" => data <= x"28";
            when "11" & x"add" => data <= x"08";
            when "11" & x"ade" => data <= x"48";
            when "11" & x"adf" => data <= x"20";
            when "11" & x"ae0" => data <= x"63";
            when "11" & x"ae1" => data <= x"af";
            when "11" & x"ae2" => data <= x"68";
            when "11" & x"ae3" => data <= x"28";
            when "11" & x"ae4" => data <= x"08";
            when "11" & x"ae5" => data <= x"48";
            when "11" & x"ae6" => data <= x"ae";
            when "11" & x"ae7" => data <= x"5b";
            when "11" & x"ae8" => data <= x"0d";
            when "11" & x"ae9" => data <= x"20";
            when "11" & x"aea" => data <= x"0f";
            when "11" & x"aeb" => data <= x"b0";
            when "11" & x"aec" => data <= x"20";
            when "11" & x"aed" => data <= x"44";
            when "11" & x"aee" => data <= x"b6";
            when "11" & x"aef" => data <= x"44";
            when "11" & x"af0" => data <= x"69";
            when "11" & x"af1" => data <= x"73";
            when "11" & x"af2" => data <= x"6b";
            when "11" & x"af3" => data <= x"20";
            when "11" & x"af4" => data <= x"00";
            when "11" & x"af5" => data <= x"68";
            when "11" & x"af6" => data <= x"28";
            when "11" & x"af7" => data <= x"20";
            when "11" & x"af8" => data <= x"6c";
            when "11" & x"af9" => data <= x"ad";
            when "11" & x"afa" => data <= x"8e";
            when "11" & x"afb" => data <= x"55";
            when "11" & x"afc" => data <= x"0d";
            when "11" & x"afd" => data <= x"a2";
            when "11" & x"afe" => data <= x"00";
            when "11" & x"aff" => data <= x"a0";
            when "11" & x"b00" => data <= x"04";
            when "11" & x"b01" => data <= x"20";
            when "11" & x"b02" => data <= x"26";
            when "11" & x"b03" => data <= x"b6";
            when "11" & x"b04" => data <= x"ad";
            when "11" & x"b05" => data <= x"55";
            when "11" & x"b06" => data <= x"0d";
            when "11" & x"b07" => data <= x"20";
            when "11" & x"b08" => data <= x"26";
            when "11" & x"b09" => data <= x"b6";
            when "11" & x"b0a" => data <= x"20";
            when "11" & x"b0b" => data <= x"44";
            when "11" & x"b0c" => data <= x"b6";
            when "11" & x"b0d" => data <= x"20";
            when "11" & x"b0e" => data <= x"69";
            when "11" & x"b0f" => data <= x"6e";
            when "11" & x"b10" => data <= x"20";
            when "11" & x"b11" => data <= x"64";
            when "11" & x"b12" => data <= x"72";
            when "11" & x"b13" => data <= x"69";
            when "11" & x"b14" => data <= x"76";
            when "11" & x"b15" => data <= x"65";
            when "11" & x"b16" => data <= x"20";
            when "11" & x"b17" => data <= x"00";
            when "11" & x"b18" => data <= x"ad";
            when "11" & x"b19" => data <= x"5b";
            when "11" & x"b1a" => data <= x"0d";
            when "11" & x"b1b" => data <= x"a2";
            when "11" & x"b1c" => data <= x"00";
            when "11" & x"b1d" => data <= x"a0";
            when "11" & x"b1e" => data <= x"02";
            when "11" & x"b1f" => data <= x"20";
            when "11" & x"b20" => data <= x"26";
            when "11" & x"b21" => data <= x"b6";
            when "11" & x"b22" => data <= x"4c";
            when "11" & x"b23" => data <= x"e7";
            when "11" & x"b24" => data <= x"ff";
            when "11" & x"b25" => data <= x"a9";
            when "11" & x"b26" => data <= x"10";
            when "11" & x"b27" => data <= x"85";
            when "11" & x"b28" => data <= x"f2";
            when "11" & x"b29" => data <= x"a9";
            when "11" & x"b2a" => data <= x"0e";
            when "11" & x"b2b" => data <= x"85";
            when "11" & x"b2c" => data <= x"f3";
            when "11" & x"b2d" => data <= x"a9";
            when "11" & x"b2e" => data <= x"80";
            when "11" & x"b2f" => data <= x"8d";
            when "11" & x"b30" => data <= x"52";
            when "11" & x"b31" => data <= x"0d";
            when "11" & x"b32" => data <= x"20";
            when "11" & x"b33" => data <= x"a1";
            when "11" & x"b34" => data <= x"b0";
            when "11" & x"b35" => data <= x"a9";
            when "11" & x"b36" => data <= x"00";
            when "11" & x"b37" => data <= x"8d";
            when "11" & x"b38" => data <= x"53";
            when "11" & x"b39" => data <= x"0d";
            when "11" & x"b3a" => data <= x"8d";
            when "11" & x"b3b" => data <= x"54";
            when "11" & x"b3c" => data <= x"0d";
            when "11" & x"b3d" => data <= x"a0";
            when "11" & x"b3e" => data <= x"0f";
            when "11" & x"b3f" => data <= x"b1";
            when "11" & x"b40" => data <= x"f2";
            when "11" & x"b41" => data <= x"10";
            when "11" & x"b42" => data <= x"0c";
            when "11" & x"b43" => data <= x"c9";
            when "11" & x"b44" => data <= x"ff";
            when "11" & x"b45" => data <= x"f0";
            when "11" & x"b46" => data <= x"36";
            when "11" & x"b47" => data <= x"ad";
            when "11" & x"b48" => data <= x"54";
            when "11" & x"b49" => data <= x"0d";
            when "11" & x"b4a" => data <= x"6a";
            when "11" & x"b4b" => data <= x"ad";
            when "11" & x"b4c" => data <= x"53";
            when "11" & x"b4d" => data <= x"0d";
            when "11" & x"b4e" => data <= x"60";
            when "11" & x"b4f" => data <= x"ee";
            when "11" & x"b50" => data <= x"53";
            when "11" & x"b51" => data <= x"0d";
            when "11" & x"b52" => data <= x"d0";
            when "11" & x"b53" => data <= x"03";
            when "11" & x"b54" => data <= x"ee";
            when "11" & x"b55" => data <= x"54";
            when "11" & x"b56" => data <= x"0d";
            when "11" & x"b57" => data <= x"18";
            when "11" & x"b58" => data <= x"a5";
            when "11" & x"b59" => data <= x"f2";
            when "11" & x"b5a" => data <= x"69";
            when "11" & x"b5b" => data <= x"10";
            when "11" & x"b5c" => data <= x"85";
            when "11" & x"b5d" => data <= x"f2";
            when "11" & x"b5e" => data <= x"d0";
            when "11" & x"b5f" => data <= x"df";
            when "11" & x"b60" => data <= x"a5";
            when "11" & x"b61" => data <= x"f3";
            when "11" & x"b62" => data <= x"49";
            when "11" & x"b63" => data <= x"01";
            when "11" & x"b64" => data <= x"85";
            when "11" & x"b65" => data <= x"f3";
            when "11" & x"b66" => data <= x"29";
            when "11" & x"b67" => data <= x"01";
            when "11" & x"b68" => data <= x"d0";
            when "11" & x"b69" => data <= x"d5";
            when "11" & x"b6a" => data <= x"18";
            when "11" & x"b6b" => data <= x"ad";
            when "11" & x"b6c" => data <= x"52";
            when "11" & x"b6d" => data <= x"0d";
            when "11" & x"b6e" => data <= x"69";
            when "11" & x"b6f" => data <= x"01";
            when "11" & x"b70" => data <= x"c9";
            when "11" & x"b71" => data <= x"90";
            when "11" & x"b72" => data <= x"f0";
            when "11" & x"b73" => data <= x"09";
            when "11" & x"b74" => data <= x"8d";
            when "11" & x"b75" => data <= x"52";
            when "11" & x"b76" => data <= x"0d";
            when "11" & x"b77" => data <= x"20";
            when "11" & x"b78" => data <= x"a1";
            when "11" & x"b79" => data <= x"b0";
            when "11" & x"b7a" => data <= x"4c";
            when "11" & x"b7b" => data <= x"3d";
            when "11" & x"b7c" => data <= x"bb";
            when "11" & x"b7d" => data <= x"20";
            when "11" & x"b7e" => data <= x"00";
            when "11" & x"b7f" => data <= x"a0";
            when "11" & x"b80" => data <= x"ff";
            when "11" & x"b81" => data <= x"4e";
            when "11" & x"b82" => data <= x"6f";
            when "11" & x"b83" => data <= x"20";
            when "11" & x"b84" => data <= x"66";
            when "11" & x"b85" => data <= x"72";
            when "11" & x"b86" => data <= x"65";
            when "11" & x"b87" => data <= x"65";
            when "11" & x"b88" => data <= x"20";
            when "11" & x"b89" => data <= x"64";
            when "11" & x"b8a" => data <= x"69";
            when "11" & x"b8b" => data <= x"73";
            when "11" & x"b8c" => data <= x"6b";
            when "11" & x"b8d" => data <= x"73";
            when "11" & x"b8e" => data <= x"00";
            when "11" & x"b8f" => data <= x"20";
            when "11" & x"b90" => data <= x"8a";
            when "11" & x"b91" => data <= x"b7";
            when "11" & x"b92" => data <= x"08";
            when "11" & x"b93" => data <= x"48";
            when "11" & x"b94" => data <= x"8a";
            when "11" & x"b95" => data <= x"48";
            when "11" & x"b96" => data <= x"a9";
            when "11" & x"b97" => data <= x"80";
            when "11" & x"b98" => data <= x"20";
            when "11" & x"b99" => data <= x"a1";
            when "11" & x"b9a" => data <= x"b0";
            when "11" & x"b9b" => data <= x"68";
            when "11" & x"b9c" => data <= x"aa";
            when "11" & x"b9d" => data <= x"68";
            when "11" & x"b9e" => data <= x"9d";
            when "11" & x"b9f" => data <= x"00";
            when "11" & x"ba0" => data <= x"0e";
            when "11" & x"ba1" => data <= x"68";
            when "11" & x"ba2" => data <= x"29";
            when "11" & x"ba3" => data <= x"01";
            when "11" & x"ba4" => data <= x"9d";
            when "11" & x"ba5" => data <= x"04";
            when "11" & x"ba6" => data <= x"0e";
            when "11" & x"ba7" => data <= x"4c";
            when "11" & x"ba8" => data <= x"b8";
            when "11" & x"ba9" => data <= x"b0";
            when "11" & x"baa" => data <= x"20";
            when "11" & x"bab" => data <= x"e4";
            when "11" & x"bac" => data <= x"bb";
            when "11" & x"bad" => data <= x"20";
            when "11" & x"bae" => data <= x"b0";
            when "11" & x"baf" => data <= x"b4";
            when "11" & x"bb0" => data <= x"a2";
            when "11" & x"bb1" => data <= x"00";
            when "11" & x"bb2" => data <= x"b0";
            when "11" & x"bb3" => data <= x"10";
            when "11" & x"bb4" => data <= x"20";
            when "11" & x"bb5" => data <= x"c3";
            when "11" & x"bb6" => data <= x"b4";
            when "11" & x"bb7" => data <= x"b0";
            when "11" & x"bb8" => data <= x"17";
            when "11" & x"bb9" => data <= x"c9";
            when "11" & x"bba" => data <= x"00";
            when "11" & x"bbb" => data <= x"d0";
            when "11" & x"bbc" => data <= x"04";
            when "11" & x"bbd" => data <= x"e0";
            when "11" & x"bbe" => data <= x"00";
            when "11" & x"bbf" => data <= x"f0";
            when "11" & x"bc0" => data <= x"03";
            when "11" & x"bc1" => data <= x"20";
            when "11" & x"bc2" => data <= x"ef";
            when "11" & x"bc3" => data <= x"bb";
            when "11" & x"bc4" => data <= x"20";
            when "11" & x"bc5" => data <= x"e2";
            when "11" & x"bc6" => data <= x"8d";
            when "11" & x"bc7" => data <= x"a2";
            when "11" & x"bc8" => data <= x"ff";
            when "11" & x"bc9" => data <= x"8a";
            when "11" & x"bca" => data <= x"8d";
            when "11" & x"bcb" => data <= x"52";
            when "11" & x"bcc" => data <= x"0d";
            when "11" & x"bcd" => data <= x"4c";
            when "11" & x"bce" => data <= x"3a";
            when "11" & x"bcf" => data <= x"b1";
            when "11" & x"bd0" => data <= x"20";
            when "11" & x"bd1" => data <= x"00";
            when "11" & x"bd2" => data <= x"a0";
            when "11" & x"bd3" => data <= x"ff";
            when "11" & x"bd4" => data <= x"42";
            when "11" & x"bd5" => data <= x"61";
            when "11" & x"bd6" => data <= x"64";
            when "11" & x"bd7" => data <= x"20";
            when "11" & x"bd8" => data <= x"66";
            when "11" & x"bd9" => data <= x"69";
            when "11" & x"bda" => data <= x"6c";
            when "11" & x"bdb" => data <= x"65";
            when "11" & x"bdc" => data <= x"20";
            when "11" & x"bdd" => data <= x"6e";
            when "11" & x"bde" => data <= x"75";
            when "11" & x"bdf" => data <= x"6d";
            when "11" & x"be0" => data <= x"62";
            when "11" & x"be1" => data <= x"65";
            when "11" & x"be2" => data <= x"72";
            when "11" & x"be3" => data <= x"00";
            when "11" & x"be4" => data <= x"a2";
            when "11" & x"be5" => data <= x"03";
            when "11" & x"be6" => data <= x"a9";
            when "11" & x"be7" => data <= x"20";
            when "11" & x"be8" => data <= x"9d";
            when "11" & x"be9" => data <= x"74";
            when "11" & x"bea" => data <= x"0d";
            when "11" & x"beb" => data <= x"ca";
            when "11" & x"bec" => data <= x"10";
            when "11" & x"bed" => data <= x"f8";
            when "11" & x"bee" => data <= x"60";
            when "11" & x"bef" => data <= x"c0";
            when "11" & x"bf0" => data <= x"09";
            when "11" & x"bf1" => data <= x"b0";
            when "11" & x"bf2" => data <= x"dd";
            when "11" & x"bf3" => data <= x"a0";
            when "11" & x"bf4" => data <= x"03";
            when "11" & x"bf5" => data <= x"b1";
            when "11" & x"bf6" => data <= x"f2";
            when "11" & x"bf7" => data <= x"29";
            when "11" & x"bf8" => data <= x"4f";
            when "11" & x"bf9" => data <= x"c9";
            when "11" & x"bfa" => data <= x"42";
            when "11" & x"bfb" => data <= x"d0";
            when "11" & x"bfc" => data <= x"d3";
            when "11" & x"bfd" => data <= x"a2";
            when "11" & x"bfe" => data <= x"00";
            when "11" & x"bff" => data <= x"c8";
            when "11" & x"c00" => data <= x"b1";
            when "11" & x"c01" => data <= x"f2";
            when "11" & x"c02" => data <= x"c9";
            when "11" & x"c03" => data <= x"20";
            when "11" & x"c04" => data <= x"f0";
            when "11" & x"c05" => data <= x"f9";
            when "11" & x"c06" => data <= x"c9";
            when "11" & x"c07" => data <= x"0d";
            when "11" & x"c08" => data <= x"f0";
            when "11" & x"c09" => data <= x"08";
            when "11" & x"c0a" => data <= x"9d";
            when "11" & x"c0b" => data <= x"74";
            when "11" & x"c0c" => data <= x"0d";
            when "11" & x"c0d" => data <= x"e8";
            when "11" & x"c0e" => data <= x"e0";
            when "11" & x"c0f" => data <= x"04";
            when "11" & x"c10" => data <= x"90";
            when "11" & x"c11" => data <= x"ed";
            when "11" & x"c12" => data <= x"a2";
            when "11" & x"c13" => data <= x"00";
            when "11" & x"c14" => data <= x"60";
            when "11" & x"c15" => data <= x"4c";
            when "11" & x"c16" => data <= x"1e";
            when "11" & x"c17" => data <= x"bc";
            when "11" & x"c18" => data <= x"4c";
            when "11" & x"c19" => data <= x"2b";
            when "11" & x"c1a" => data <= x"bc";
            when "11" & x"c1b" => data <= x"4c";
            when "11" & x"c1c" => data <= x"38";
            when "11" & x"c1d" => data <= x"bc";
            when "11" & x"c1e" => data <= x"20";
            when "11" & x"c1f" => data <= x"d8";
            when "11" & x"c20" => data <= x"bd";
            when "11" & x"c21" => data <= x"20";
            when "11" & x"c22" => data <= x"a7";
            when "11" & x"c23" => data <= x"bd";
            when "11" & x"c24" => data <= x"20";
            when "11" & x"c25" => data <= x"d0";
            when "11" & x"c26" => data <= x"bd";
            when "11" & x"c27" => data <= x"20";
            when "11" & x"c28" => data <= x"05";
            when "11" & x"c29" => data <= x"be";
            when "11" & x"c2a" => data <= x"60";
            when "11" & x"c2b" => data <= x"20";
            when "11" & x"c2c" => data <= x"d8";
            when "11" & x"c2d" => data <= x"bd";
            when "11" & x"c2e" => data <= x"20";
            when "11" & x"c2f" => data <= x"a7";
            when "11" & x"c30" => data <= x"bd";
            when "11" & x"c31" => data <= x"20";
            when "11" & x"c32" => data <= x"d4";
            when "11" & x"c33" => data <= x"bd";
            when "11" & x"c34" => data <= x"20";
            when "11" & x"c35" => data <= x"05";
            when "11" & x"c36" => data <= x"be";
            when "11" & x"c37" => data <= x"60";
            when "11" & x"c38" => data <= x"a9";
            when "11" & x"c39" => data <= x"00";
            when "11" & x"c3a" => data <= x"8d";
            when "11" & x"c3b" => data <= x"28";
            when "11" & x"c3c" => data <= x"0d";
            when "11" & x"c3d" => data <= x"20";
            when "11" & x"c3e" => data <= x"c2";
            when "11" & x"c3f" => data <= x"ff";
            when "11" & x"c40" => data <= x"f0";
            when "11" & x"c41" => data <= x"6e";
            when "11" & x"c42" => data <= x"b1";
            when "11" & x"c43" => data <= x"f2";
            when "11" & x"c44" => data <= x"c8";
            when "11" & x"c45" => data <= x"c9";
            when "11" & x"c46" => data <= x"20";
            when "11" & x"c47" => data <= x"f0";
            when "11" & x"c48" => data <= x"f9";
            when "11" & x"c49" => data <= x"b1";
            when "11" & x"c4a" => data <= x"f2";
            when "11" & x"c4b" => data <= x"88";
            when "11" & x"c4c" => data <= x"c9";
            when "11" & x"c4d" => data <= x"20";
            when "11" & x"c4e" => data <= x"d0";
            when "11" & x"c4f" => data <= x"24";
            when "11" & x"c50" => data <= x"b1";
            when "11" & x"c51" => data <= x"f2";
            when "11" & x"c52" => data <= x"38";
            when "11" & x"c53" => data <= x"e9";
            when "11" & x"c54" => data <= x"30";
            when "11" & x"c55" => data <= x"30";
            when "11" & x"c56" => data <= x"1d";
            when "11" & x"c57" => data <= x"c9";
            when "11" & x"c58" => data <= x"0a";
            when "11" & x"c59" => data <= x"90";
            when "11" & x"c5a" => data <= x"14";
            when "11" & x"c5b" => data <= x"e9";
            when "11" & x"c5c" => data <= x"07";
            when "11" & x"c5d" => data <= x"c9";
            when "11" & x"c5e" => data <= x"0a";
            when "11" & x"c5f" => data <= x"90";
            when "11" & x"c60" => data <= x"13";
            when "11" & x"c61" => data <= x"c9";
            when "11" & x"c62" => data <= x"10";
            when "11" & x"c63" => data <= x"90";
            when "11" & x"c64" => data <= x"0a";
            when "11" & x"c65" => data <= x"e9";
            when "11" & x"c66" => data <= x"20";
            when "11" & x"c67" => data <= x"c9";
            when "11" & x"c68" => data <= x"0a";
            when "11" & x"c69" => data <= x"90";
            when "11" & x"c6a" => data <= x"09";
            when "11" & x"c6b" => data <= x"c9";
            when "11" & x"c6c" => data <= x"10";
            when "11" & x"c6d" => data <= x"b0";
            when "11" & x"c6e" => data <= x"05";
            when "11" & x"c6f" => data <= x"c8";
            when "11" & x"c70" => data <= x"c8";
            when "11" & x"c71" => data <= x"8d";
            when "11" & x"c72" => data <= x"28";
            when "11" & x"c73" => data <= x"0d";
            when "11" & x"c74" => data <= x"a5";
            when "11" & x"c75" => data <= x"f4";
            when "11" & x"c76" => data <= x"8d";
            when "11" & x"c77" => data <= x"29";
            when "11" & x"c78" => data <= x"0d";
            when "11" & x"c79" => data <= x"98";
            when "11" & x"c7a" => data <= x"48";
            when "11" & x"c7b" => data <= x"a0";
            when "11" & x"c7c" => data <= x"26";
            when "11" & x"c7d" => data <= x"b9";
            when "11" & x"c7e" => data <= x"81";
            when "11" & x"c7f" => data <= x"bd";
            when "11" & x"c80" => data <= x"99";
            when "11" & x"c81" => data <= x"52";
            when "11" & x"c82" => data <= x"0d";
            when "11" & x"c83" => data <= x"88";
            when "11" & x"c84" => data <= x"10";
            when "11" & x"c85" => data <= x"f7";
            when "11" & x"c86" => data <= x"a2";
            when "11" & x"c87" => data <= x"0f";
            when "11" & x"c88" => data <= x"20";
            when "11" & x"c89" => data <= x"52";
            when "11" & x"c8a" => data <= x"0d";
            when "11" & x"c8b" => data <= x"68";
            when "11" & x"c8c" => data <= x"a8";
            when "11" & x"c8d" => data <= x"8e";
            when "11" & x"c8e" => data <= x"28";
            when "11" & x"c8f" => data <= x"0d";
            when "11" & x"c90" => data <= x"8a";
            when "11" & x"c91" => data <= x"10";
            when "11" & x"c92" => data <= x"14";
            when "11" & x"c93" => data <= x"20";
            when "11" & x"c94" => data <= x"00";
            when "11" & x"c95" => data <= x"a0";
            when "11" & x"c96" => data <= x"ff";
            when "11" & x"c97" => data <= x"4e";
            when "11" & x"c98" => data <= x"6f";
            when "11" & x"c99" => data <= x"20";
            when "11" & x"c9a" => data <= x"53";
            when "11" & x"c9b" => data <= x"69";
            when "11" & x"c9c" => data <= x"64";
            when "11" & x"c9d" => data <= x"65";
            when "11" & x"c9e" => data <= x"77";
            when "11" & x"c9f" => data <= x"61";
            when "11" & x"ca0" => data <= x"79";
            when "11" & x"ca1" => data <= x"73";
            when "11" & x"ca2" => data <= x"20";
            when "11" & x"ca3" => data <= x"52";
            when "11" & x"ca4" => data <= x"41";
            when "11" & x"ca5" => data <= x"4d";
            when "11" & x"ca6" => data <= x"00";
            when "11" & x"ca7" => data <= x"20";
            when "11" & x"ca8" => data <= x"62";
            when "11" & x"ca9" => data <= x"82";
            when "11" & x"caa" => data <= x"18";
            when "11" & x"cab" => data <= x"20";
            when "11" & x"cac" => data <= x"c2";
            when "11" & x"cad" => data <= x"ff";
            when "11" & x"cae" => data <= x"d0";
            when "11" & x"caf" => data <= x"03";
            when "11" & x"cb0" => data <= x"4c";
            when "11" & x"cb1" => data <= x"f5";
            when "11" & x"cb2" => data <= x"b6";
            when "11" & x"cb3" => data <= x"20";
            when "11" & x"cb4" => data <= x"fe";
            when "11" & x"cb5" => data <= x"80";
            when "11" & x"cb6" => data <= x"98";
            when "11" & x"cb7" => data <= x"20";
            when "11" & x"cb8" => data <= x"71";
            when "11" & x"cb9" => data <= x"82";
            when "11" & x"cba" => data <= x"b9";
            when "11" & x"cbb" => data <= x"0e";
            when "11" & x"cbc" => data <= x"0f";
            when "11" & x"cbd" => data <= x"48";
            when "11" & x"cbe" => data <= x"29";
            when "11" & x"cbf" => data <= x"03";
            when "11" & x"cc0" => data <= x"85";
            when "11" & x"cc1" => data <= x"a1";
            when "11" & x"cc2" => data <= x"b9";
            when "11" & x"cc3" => data <= x"0f";
            when "11" & x"cc4" => data <= x"0f";
            when "11" & x"cc5" => data <= x"85";
            when "11" & x"cc6" => data <= x"a0";
            when "11" & x"cc7" => data <= x"68";
            when "11" & x"cc8" => data <= x"4a";
            when "11" & x"cc9" => data <= x"4a";
            when "11" & x"cca" => data <= x"29";
            when "11" & x"ccb" => data <= x"03";
            when "11" & x"ccc" => data <= x"f0";
            when "11" & x"ccd" => data <= x"04";
            when "11" & x"cce" => data <= x"49";
            when "11" & x"ccf" => data <= x"03";
            when "11" & x"cd0" => data <= x"d0";
            when "11" & x"cd1" => data <= x"17";
            when "11" & x"cd2" => data <= x"b9";
            when "11" & x"cd3" => data <= x"0c";
            when "11" & x"cd4" => data <= x"0f";
            when "11" & x"cd5" => data <= x"d0";
            when "11" & x"cd6" => data <= x"12";
            when "11" & x"cd7" => data <= x"b9";
            when "11" & x"cd8" => data <= x"0d";
            when "11" & x"cd9" => data <= x"0f";
            when "11" & x"cda" => data <= x"30";
            when "11" & x"cdb" => data <= x"0d";
            when "11" & x"cdc" => data <= x"8d";
            when "11" & x"cdd" => data <= x"27";
            when "11" & x"cde" => data <= x"0d";
            when "11" & x"cdf" => data <= x"a2";
            when "11" & x"ce0" => data <= x"05";
            when "11" & x"ce1" => data <= x"c9";
            when "11" & x"ce2" => data <= x"40";
            when "11" & x"ce3" => data <= x"f0";
            when "11" & x"ce4" => data <= x"15";
            when "11" & x"ce5" => data <= x"0a";
            when "11" & x"ce6" => data <= x"ca";
            when "11" & x"ce7" => data <= x"d0";
            when "11" & x"ce8" => data <= x"f8";
            when "11" & x"ce9" => data <= x"20";
            when "11" & x"cea" => data <= x"00";
            when "11" & x"ceb" => data <= x"a0";
            when "11" & x"cec" => data <= x"ff";
            when "11" & x"ced" => data <= x"42";
            when "11" & x"cee" => data <= x"61";
            when "11" & x"cef" => data <= x"64";
            when "11" & x"cf0" => data <= x"20";
            when "11" & x"cf1" => data <= x"52";
            when "11" & x"cf2" => data <= x"4f";
            when "11" & x"cf3" => data <= x"4d";
            when "11" & x"cf4" => data <= x"20";
            when "11" & x"cf5" => data <= x"73";
            when "11" & x"cf6" => data <= x"69";
            when "11" & x"cf7" => data <= x"7a";
            when "11" & x"cf8" => data <= x"65";
            when "11" & x"cf9" => data <= x"00";
            when "11" & x"cfa" => data <= x"4e";
            when "11" & x"cfb" => data <= x"27";
            when "11" & x"cfc" => data <= x"0d";
            when "11" & x"cfd" => data <= x"a6";
            when "11" & x"cfe" => data <= x"cf";
            when "11" & x"cff" => data <= x"20";
            when "11" & x"d00" => data <= x"1d";
            when "11" & x"d01" => data <= x"ae";
            when "11" & x"d02" => data <= x"18";
            when "11" & x"d03" => data <= x"ad";
            when "11" & x"d04" => data <= x"23";
            when "11" & x"d05" => data <= x"0d";
            when "11" & x"d06" => data <= x"65";
            when "11" & x"d07" => data <= x"a0";
            when "11" & x"d08" => data <= x"8d";
            when "11" & x"d09" => data <= x"23";
            when "11" & x"d0a" => data <= x"0d";
            when "11" & x"d0b" => data <= x"ad";
            when "11" & x"d0c" => data <= x"24";
            when "11" & x"d0d" => data <= x"0d";
            when "11" & x"d0e" => data <= x"65";
            when "11" & x"d0f" => data <= x"a1";
            when "11" & x"d10" => data <= x"8d";
            when "11" & x"d11" => data <= x"24";
            when "11" & x"d12" => data <= x"0d";
            when "11" & x"d13" => data <= x"a9";
            when "11" & x"d14" => data <= x"00";
            when "11" & x"d15" => data <= x"6d";
            when "11" & x"d16" => data <= x"25";
            when "11" & x"d17" => data <= x"0d";
            when "11" & x"d18" => data <= x"8d";
            when "11" & x"d19" => data <= x"25";
            when "11" & x"d1a" => data <= x"0d";
            when "11" & x"d1b" => data <= x"a0";
            when "11" & x"d1c" => data <= x"1c";
            when "11" & x"d1d" => data <= x"b9";
            when "11" & x"d1e" => data <= x"65";
            when "11" & x"d1f" => data <= x"bd";
            when "11" & x"d20" => data <= x"99";
            when "11" & x"d21" => data <= x"52";
            when "11" & x"d22" => data <= x"0d";
            when "11" & x"d23" => data <= x"88";
            when "11" & x"d24" => data <= x"10";
            when "11" & x"d25" => data <= x"f7";
            when "11" & x"d26" => data <= x"ad";
            when "11" & x"d27" => data <= x"28";
            when "11" & x"d28" => data <= x"0d";
            when "11" & x"d29" => data <= x"8d";
            when "11" & x"d2a" => data <= x"53";
            when "11" & x"d2b" => data <= x"0d";
            when "11" & x"d2c" => data <= x"ad";
            when "11" & x"d2d" => data <= x"29";
            when "11" & x"d2e" => data <= x"0d";
            when "11" & x"d2f" => data <= x"8d";
            when "11" & x"d30" => data <= x"69";
            when "11" & x"d31" => data <= x"0d";
            when "11" & x"d32" => data <= x"20";
            when "11" & x"d33" => data <= x"1f";
            when "11" & x"d34" => data <= x"a6";
            when "11" & x"d35" => data <= x"a9";
            when "11" & x"d36" => data <= x"ff";
            when "11" & x"d37" => data <= x"8d";
            when "11" & x"d38" => data <= x"82";
            when "11" & x"d39" => data <= x"10";
            when "11" & x"d3a" => data <= x"20";
            when "11" & x"d3b" => data <= x"99";
            when "11" & x"d3c" => data <= x"a7";
            when "11" & x"d3d" => data <= x"20";
            when "11" & x"d3e" => data <= x"52";
            when "11" & x"d3f" => data <= x"0d";
            when "11" & x"d40" => data <= x"18";
            when "11" & x"d41" => data <= x"ad";
            when "11" & x"d42" => data <= x"23";
            when "11" & x"d43" => data <= x"0d";
            when "11" & x"d44" => data <= x"69";
            when "11" & x"d45" => data <= x"02";
            when "11" & x"d46" => data <= x"8d";
            when "11" & x"d47" => data <= x"23";
            when "11" & x"d48" => data <= x"0d";
            when "11" & x"d49" => data <= x"90";
            when "11" & x"d4a" => data <= x"08";
            when "11" & x"d4b" => data <= x"ee";
            when "11" & x"d4c" => data <= x"24";
            when "11" & x"d4d" => data <= x"0d";
            when "11" & x"d4e" => data <= x"d0";
            when "11" & x"d4f" => data <= x"03";
            when "11" & x"d50" => data <= x"ee";
            when "11" & x"d51" => data <= x"24";
            when "11" & x"d52" => data <= x"0d";
            when "11" & x"d53" => data <= x"ee";
            when "11" & x"d54" => data <= x"5e";
            when "11" & x"d55" => data <= x"0d";
            when "11" & x"d56" => data <= x"ee";
            when "11" & x"d57" => data <= x"5e";
            when "11" & x"d58" => data <= x"0d";
            when "11" & x"d59" => data <= x"ee";
            when "11" & x"d5a" => data <= x"64";
            when "11" & x"d5b" => data <= x"0d";
            when "11" & x"d5c" => data <= x"ee";
            when "11" & x"d5d" => data <= x"64";
            when "11" & x"d5e" => data <= x"0d";
            when "11" & x"d5f" => data <= x"ce";
            when "11" & x"d60" => data <= x"27";
            when "11" & x"d61" => data <= x"0d";
            when "11" & x"d62" => data <= x"d0";
            when "11" & x"d63" => data <= x"d6";
            when "11" & x"d64" => data <= x"60";
            when "11" & x"d65" => data <= x"a9";
            when "11" & x"d66" => data <= x"00";
            when "11" & x"d67" => data <= x"8d";
            when "11" & x"d68" => data <= x"30";
            when "11" & x"d69" => data <= x"fe";
            when "11" & x"d6a" => data <= x"a0";
            when "11" & x"d6b" => data <= x"00";
            when "11" & x"d6c" => data <= x"b9";
            when "11" & x"d6d" => data <= x"00";
            when "11" & x"d6e" => data <= x"0e";
            when "11" & x"d6f" => data <= x"99";
            when "11" & x"d70" => data <= x"00";
            when "11" & x"d71" => data <= x"80";
            when "11" & x"d72" => data <= x"b9";
            when "11" & x"d73" => data <= x"00";
            when "11" & x"d74" => data <= x"0f";
            when "11" & x"d75" => data <= x"99";
            when "11" & x"d76" => data <= x"00";
            when "11" & x"d77" => data <= x"81";
            when "11" & x"d78" => data <= x"88";
            when "11" & x"d79" => data <= x"d0";
            when "11" & x"d7a" => data <= x"f1";
            when "11" & x"d7b" => data <= x"a9";
            when "11" & x"d7c" => data <= x"00";
            when "11" & x"d7d" => data <= x"8d";
            when "11" & x"d7e" => data <= x"30";
            when "11" & x"d7f" => data <= x"fe";
            when "11" & x"d80" => data <= x"60";
            when "11" & x"d81" => data <= x"8e";
            when "11" & x"d82" => data <= x"30";
            when "11" & x"d83" => data <= x"fe";
            when "11" & x"d84" => data <= x"ad";
            when "11" & x"d85" => data <= x"ff";
            when "11" & x"d86" => data <= x"bf";
            when "11" & x"d87" => data <= x"a8";
            when "11" & x"d88" => data <= x"49";
            when "11" & x"d89" => data <= x"ff";
            when "11" & x"d8a" => data <= x"8d";
            when "11" & x"d8b" => data <= x"ff";
            when "11" & x"d8c" => data <= x"bf";
            when "11" & x"d8d" => data <= x"98";
            when "11" & x"d8e" => data <= x"4d";
            when "11" & x"d8f" => data <= x"ff";
            when "11" & x"d90" => data <= x"bf";
            when "11" & x"d91" => data <= x"8c";
            when "11" & x"d92" => data <= x"ff";
            when "11" & x"d93" => data <= x"bf";
            when "11" & x"d94" => data <= x"c9";
            when "11" & x"d95" => data <= x"ff";
            when "11" & x"d96" => data <= x"d0";
            when "11" & x"d97" => data <= x"05";
            when "11" & x"d98" => data <= x"ce";
            when "11" & x"d99" => data <= x"28";
            when "11" & x"d9a" => data <= x"0d";
            when "11" & x"d9b" => data <= x"30";
            when "11" & x"d9c" => data <= x"03";
            when "11" & x"d9d" => data <= x"ca";
            when "11" & x"d9e" => data <= x"10";
            when "11" & x"d9f" => data <= x"e1";
            when "11" & x"da0" => data <= x"ad";
            when "11" & x"da1" => data <= x"29";
            when "11" & x"da2" => data <= x"0d";
            when "11" & x"da3" => data <= x"8d";
            when "11" & x"da4" => data <= x"30";
            when "11" & x"da5" => data <= x"fe";
            when "11" & x"da6" => data <= x"60";
            when "11" & x"da7" => data <= x"a2";
            when "11" & x"da8" => data <= x"0b";
            when "11" & x"da9" => data <= x"bd";
            when "11" & x"daa" => data <= x"32";
            when "11" & x"dab" => data <= x"be";
            when "11" & x"dac" => data <= x"9d";
            when "11" & x"dad" => data <= x"70";
            when "11" & x"dae" => data <= x"0d";
            when "11" & x"daf" => data <= x"ca";
            when "11" & x"db0" => data <= x"10";
            when "11" & x"db1" => data <= x"f7";
            when "11" & x"db2" => data <= x"e8";
            when "11" & x"db3" => data <= x"8e";
            when "11" & x"db4" => data <= x"05";
            when "11" & x"db5" => data <= x"0d";
            when "11" & x"db6" => data <= x"8e";
            when "11" & x"db7" => data <= x"28";
            when "11" & x"db8" => data <= x"0d";
            when "11" & x"db9" => data <= x"a9";
            when "11" & x"dba" => data <= x"40";
            when "11" & x"dbb" => data <= x"8d";
            when "11" & x"dbc" => data <= x"27";
            when "11" & x"dbd" => data <= x"0d";
            when "11" & x"dbe" => data <= x"0a";
            when "11" & x"dbf" => data <= x"48";
            when "11" & x"dc0" => data <= x"20";
            when "11" & x"dc1" => data <= x"1f";
            when "11" & x"dc2" => data <= x"a6";
            when "11" & x"dc3" => data <= x"68";
            when "11" & x"dc4" => data <= x"20";
            when "11" & x"dc5" => data <= x"70";
            when "11" & x"dc6" => data <= x"b0";
            when "11" & x"dc7" => data <= x"a9";
            when "11" & x"dc8" => data <= x"00";
            when "11" & x"dc9" => data <= x"85";
            when "11" & x"dca" => data <= x"a0";
            when "11" & x"dcb" => data <= x"a9";
            when "11" & x"dcc" => data <= x"20";
            when "11" & x"dcd" => data <= x"85";
            when "11" & x"dce" => data <= x"a1";
            when "11" & x"dcf" => data <= x"60";
            when "11" & x"dd0" => data <= x"20";
            when "11" & x"dd1" => data <= x"cc";
            when "11" & x"dd2" => data <= x"a7";
            when "11" & x"dd3" => data <= x"60";
            when "11" & x"dd4" => data <= x"20";
            when "11" & x"dd5" => data <= x"78";
            when "11" & x"dd6" => data <= x"a8";
            when "11" & x"dd7" => data <= x"60";
            when "11" & x"dd8" => data <= x"a2";
            when "11" & x"dd9" => data <= x"0b";
            when "11" & x"dda" => data <= x"bd";
            when "11" & x"ddb" => data <= x"70";
            when "11" & x"ddc" => data <= x"0d";
            when "11" & x"ddd" => data <= x"9d";
            when "11" & x"dde" => data <= x"60";
            when "11" & x"ddf" => data <= x"0d";
            when "11" & x"de0" => data <= x"ca";
            when "11" & x"de1" => data <= x"10";
            when "11" & x"de2" => data <= x"f7";
            when "11" & x"de3" => data <= x"a2";
            when "11" & x"de4" => data <= x"06";
            when "11" & x"de5" => data <= x"bd";
            when "11" & x"de6" => data <= x"05";
            when "11" & x"de7" => data <= x"0d";
            when "11" & x"de8" => data <= x"9d";
            when "11" & x"de9" => data <= x"2e";
            when "11" & x"dea" => data <= x"0d";
            when "11" & x"deb" => data <= x"ca";
            when "11" & x"dec" => data <= x"10";
            when "11" & x"ded" => data <= x"f7";
            when "11" & x"dee" => data <= x"ad";
            when "11" & x"def" => data <= x"28";
            when "11" & x"df0" => data <= x"0d";
            when "11" & x"df1" => data <= x"8d";
            when "11" & x"df2" => data <= x"35";
            when "11" & x"df3" => data <= x"0d";
            when "11" & x"df4" => data <= x"a5";
            when "11" & x"df5" => data <= x"a0";
            when "11" & x"df6" => data <= x"8d";
            when "11" & x"df7" => data <= x"36";
            when "11" & x"df8" => data <= x"0d";
            when "11" & x"df9" => data <= x"a5";
            when "11" & x"dfa" => data <= x"a1";
            when "11" & x"dfb" => data <= x"8d";
            when "11" & x"dfc" => data <= x"37";
            when "11" & x"dfd" => data <= x"0d";
            when "11" & x"dfe" => data <= x"ad";
            when "11" & x"dff" => data <= x"27";
            when "11" & x"e00" => data <= x"0d";
            when "11" & x"e01" => data <= x"8d";
            when "11" & x"e02" => data <= x"38";
            when "11" & x"e03" => data <= x"0d";
            when "11" & x"e04" => data <= x"60";
            when "11" & x"e05" => data <= x"ad";
            when "11" & x"e06" => data <= x"38";
            when "11" & x"e07" => data <= x"0d";
            when "11" & x"e08" => data <= x"8d";
            when "11" & x"e09" => data <= x"27";
            when "11" & x"e0a" => data <= x"0d";
            when "11" & x"e0b" => data <= x"ad";
            when "11" & x"e0c" => data <= x"37";
            when "11" & x"e0d" => data <= x"0d";
            when "11" & x"e0e" => data <= x"85";
            when "11" & x"e0f" => data <= x"a1";
            when "11" & x"e10" => data <= x"ad";
            when "11" & x"e11" => data <= x"36";
            when "11" & x"e12" => data <= x"0d";
            when "11" & x"e13" => data <= x"85";
            when "11" & x"e14" => data <= x"a0";
            when "11" & x"e15" => data <= x"ad";
            when "11" & x"e16" => data <= x"35";
            when "11" & x"e17" => data <= x"0d";
            when "11" & x"e18" => data <= x"8d";
            when "11" & x"e19" => data <= x"28";
            when "11" & x"e1a" => data <= x"0d";
            when "11" & x"e1b" => data <= x"a2";
            when "11" & x"e1c" => data <= x"06";
            when "11" & x"e1d" => data <= x"bd";
            when "11" & x"e1e" => data <= x"2e";
            when "11" & x"e1f" => data <= x"0d";
            when "11" & x"e20" => data <= x"9d";
            when "11" & x"e21" => data <= x"05";
            when "11" & x"e22" => data <= x"0d";
            when "11" & x"e23" => data <= x"ca";
            when "11" & x"e24" => data <= x"10";
            when "11" & x"e25" => data <= x"f7";
            when "11" & x"e26" => data <= x"a2";
            when "11" & x"e27" => data <= x"0b";
            when "11" & x"e28" => data <= x"bd";
            when "11" & x"e29" => data <= x"60";
            when "11" & x"e2a" => data <= x"0d";
            when "11" & x"e2b" => data <= x"9d";
            when "11" & x"e2c" => data <= x"70";
            when "11" & x"e2d" => data <= x"0d";
            when "11" & x"e2e" => data <= x"ca";
            when "11" & x"e2f" => data <= x"10";
            when "11" & x"e30" => data <= x"f7";
            when "11" & x"e31" => data <= x"60";
            when "11" & x"e32" => data <= x"49";
            when "11" & x"e33" => data <= x"4e";
            when "11" & x"e34" => data <= x"4f";
            when "11" & x"e35" => data <= x"55";
            when "11" & x"e36" => data <= x"54";
            when "11" & x"e37" => data <= x"4d";
            when "11" & x"e38" => data <= x"45";
            when "11" & x"e39" => data <= x"4d";
            when "11" & x"e3a" => data <= x"20";
            when "11" & x"e3b" => data <= x"20";
            when "11" & x"e3c" => data <= x"20";
            when "11" & x"e3d" => data <= x"20";
            when "11" & x"e3e" => data <= x"48";
            when "11" & x"e3f" => data <= x"a5";
            when "11" & x"e40" => data <= x"cf";
            when "11" & x"e41" => data <= x"8d";
            when "11" & x"e42" => data <= x"20";
            when "11" & x"e43" => data <= x"0d";
            when "11" & x"e44" => data <= x"68";
            when "11" & x"e45" => data <= x"60";
            when "11" & x"e46" => data <= x"a0";
            when "11" & x"e47" => data <= x"00";
            when "11" & x"e48" => data <= x"b1";
            when "11" & x"e49" => data <= x"b0";
            when "11" & x"e4a" => data <= x"30";
            when "11" & x"e4b" => data <= x"07";
            when "11" & x"e4c" => data <= x"29";
            when "11" & x"e4d" => data <= x"03";
            when "11" & x"e4e" => data <= x"85";
            when "11" & x"e4f" => data <= x"cf";
            when "11" & x"e50" => data <= x"8d";
            when "11" & x"e51" => data <= x"20";
            when "11" & x"e52" => data <= x"0d";
            when "11" & x"e53" => data <= x"a0";
            when "11" & x"e54" => data <= x"05";
            when "11" & x"e55" => data <= x"b1";
            when "11" & x"e56" => data <= x"b0";
            when "11" & x"e57" => data <= x"18";
            when "11" & x"e58" => data <= x"69";
            when "11" & x"e59" => data <= x"07";
            when "11" & x"e5a" => data <= x"85";
            when "11" & x"e5b" => data <= x"be";
            when "11" & x"e5c" => data <= x"20";
            when "11" & x"e5d" => data <= x"6a";
            when "11" & x"e5e" => data <= x"be";
            when "11" & x"e5f" => data <= x"a4";
            when "11" & x"e60" => data <= x"be";
            when "11" & x"e61" => data <= x"b0";
            when "11" & x"e62" => data <= x"02";
            when "11" & x"e63" => data <= x"a9";
            when "11" & x"e64" => data <= x"00";
            when "11" & x"e65" => data <= x"91";
            when "11" & x"e66" => data <= x"b0";
            when "11" & x"e67" => data <= x"a9";
            when "11" & x"e68" => data <= x"00";
            when "11" & x"e69" => data <= x"60";
            when "11" & x"e6a" => data <= x"c8";
            when "11" & x"e6b" => data <= x"b1";
            when "11" & x"e6c" => data <= x"b0";
            when "11" & x"e6d" => data <= x"aa";
            when "11" & x"e6e" => data <= x"29";
            when "11" & x"e6f" => data <= x"3f";
            when "11" & x"e70" => data <= x"85";
            when "11" & x"e71" => data <= x"bf";
            when "11" & x"e72" => data <= x"c9";
            when "11" & x"e73" => data <= x"3a";
            when "11" & x"e74" => data <= x"d0";
            when "11" & x"e75" => data <= x"2f";
            when "11" & x"e76" => data <= x"a5";
            when "11" & x"e77" => data <= x"be";
            when "11" & x"e78" => data <= x"c9";
            when "11" & x"e79" => data <= x"09";
            when "11" & x"e7a" => data <= x"d0";
            when "11" & x"e7b" => data <= x"13";
            when "11" & x"e7c" => data <= x"c8";
            when "11" & x"e7d" => data <= x"b1";
            when "11" & x"e7e" => data <= x"b0";
            when "11" & x"e7f" => data <= x"c9";
            when "11" & x"e80" => data <= x"23";
            when "11" & x"e81" => data <= x"d0";
            when "11" & x"e82" => data <= x"0c";
            when "11" & x"e83" => data <= x"c8";
            when "11" & x"e84" => data <= x"b1";
            when "11" & x"e85" => data <= x"b0";
            when "11" & x"e86" => data <= x"29";
            when "11" & x"e87" => data <= x"20";
            when "11" & x"e88" => data <= x"f0";
            when "11" & x"e89" => data <= x"02";
            when "11" & x"e8a" => data <= x"a9";
            when "11" & x"e8b" => data <= x"02";
            when "11" & x"e8c" => data <= x"8d";
            when "11" & x"e8d" => data <= x"20";
            when "11" & x"e8e" => data <= x"0d";
            when "11" & x"e8f" => data <= x"18";
            when "11" & x"e90" => data <= x"60";
            when "11" & x"e91" => data <= x"a9";
            when "11" & x"e92" => data <= x"1e";
            when "11" & x"e93" => data <= x"38";
            when "11" & x"e94" => data <= x"60";
            when "11" & x"e95" => data <= x"a9";
            when "11" & x"e96" => data <= x"10";
            when "11" & x"e97" => data <= x"38";
            when "11" & x"e98" => data <= x"60";
            when "11" & x"e99" => data <= x"a9";
            when "11" & x"e9a" => data <= x"12";
            when "11" & x"e9b" => data <= x"38";
            when "11" & x"e9c" => data <= x"60";
            when "11" & x"e9d" => data <= x"a9";
            when "11" & x"e9e" => data <= x"ff";
            when "11" & x"e9f" => data <= x"38";
            when "11" & x"ea0" => data <= x"60";
            when "11" & x"ea1" => data <= x"a9";
            when "11" & x"ea2" => data <= x"1e";
            when "11" & x"ea3" => data <= x"38";
            when "11" & x"ea4" => data <= x"60";
            when "11" & x"ea5" => data <= x"a5";
            when "11" & x"ea6" => data <= x"cf";
            when "11" & x"ea7" => data <= x"6a";
            when "11" & x"ea8" => data <= x"8a";
            when "11" & x"ea9" => data <= x"90";
            when "11" & x"eaa" => data <= x"02";
            when "11" & x"eab" => data <= x"49";
            when "11" & x"eac" => data <= x"c0";
            when "11" & x"ead" => data <= x"2a";
            when "11" & x"eae" => data <= x"90";
            when "11" & x"eaf" => data <= x"0c";
            when "11" & x"eb0" => data <= x"2a";
            when "11" & x"eb1" => data <= x"b0";
            when "11" & x"eb2" => data <= x"de";
            when "11" & x"eb3" => data <= x"ad";
            when "11" & x"eb4" => data <= x"20";
            when "11" & x"eb5" => data <= x"0d";
            when "11" & x"eb6" => data <= x"29";
            when "11" & x"eb7" => data <= x"02";
            when "11" & x"eb8" => data <= x"09";
            when "11" & x"eb9" => data <= x"01";
            when "11" & x"eba" => data <= x"d0";
            when "11" & x"ebb" => data <= x"08";
            when "11" & x"ebc" => data <= x"2a";
            when "11" & x"ebd" => data <= x"90";
            when "11" & x"ebe" => data <= x"d6";
            when "11" & x"ebf" => data <= x"ad";
            when "11" & x"ec0" => data <= x"20";
            when "11" & x"ec1" => data <= x"0d";
            when "11" & x"ec2" => data <= x"29";
            when "11" & x"ec3" => data <= x"02";
            when "11" & x"ec4" => data <= x"8d";
            when "11" & x"ec5" => data <= x"20";
            when "11" & x"ec6" => data <= x"0d";
            when "11" & x"ec7" => data <= x"aa";
            when "11" & x"ec8" => data <= x"86";
            when "11" & x"ec9" => data <= x"c0";
            when "11" & x"eca" => data <= x"bd";
            when "11" & x"ecb" => data <= x"10";
            when "11" & x"ecc" => data <= x"0d";
            when "11" & x"ecd" => data <= x"30";
            when "11" & x"ece" => data <= x"c6";
            when "11" & x"ecf" => data <= x"a5";
            when "11" & x"ed0" => data <= x"bf";
            when "11" & x"ed1" => data <= x"c9";
            when "11" & x"ed2" => data <= x"13";
            when "11" & x"ed3" => data <= x"f0";
            when "11" & x"ed4" => data <= x"0b";
            when "11" & x"ed5" => data <= x"c9";
            when "11" & x"ed6" => data <= x"0b";
            when "11" & x"ed7" => data <= x"d0";
            when "11" & x"ed8" => data <= x"b6";
            when "11" & x"ed9" => data <= x"bd";
            when "11" & x"eda" => data <= x"1c";
            when "11" & x"edb" => data <= x"0d";
            when "11" & x"edc" => data <= x"c9";
            when "11" & x"edd" => data <= x"54";
            when "11" & x"ede" => data <= x"d0";
            when "11" & x"edf" => data <= x"b9";
            when "11" & x"ee0" => data <= x"a5";
            when "11" & x"ee1" => data <= x"be";
            when "11" & x"ee2" => data <= x"c9";
            when "11" & x"ee3" => data <= x"0a";
            when "11" & x"ee4" => data <= x"d0";
            when "11" & x"ee5" => data <= x"b7";
            when "11" & x"ee6" => data <= x"20";
            when "11" & x"ee7" => data <= x"1f";
            when "11" & x"ee8" => data <= x"a6";
            when "11" & x"ee9" => data <= x"a9";
            when "11" & x"eea" => data <= x"00";
            when "11" & x"eeb" => data <= x"85";
            when "11" & x"eec" => data <= x"c5";
            when "11" & x"eed" => data <= x"c8";
            when "11" & x"eee" => data <= x"b1";
            when "11" & x"eef" => data <= x"b0";
            when "11" & x"ef0" => data <= x"c9";
            when "11" & x"ef1" => data <= x"50";
            when "11" & x"ef2" => data <= x"b0";
            when "11" & x"ef3" => data <= x"9d";
            when "11" & x"ef4" => data <= x"0a";
            when "11" & x"ef5" => data <= x"85";
            when "11" & x"ef6" => data <= x"c4";
            when "11" & x"ef7" => data <= x"0a";
            when "11" & x"ef8" => data <= x"26";
            when "11" & x"ef9" => data <= x"c5";
            when "11" & x"efa" => data <= x"0a";
            when "11" & x"efb" => data <= x"26";
            when "11" & x"efc" => data <= x"c5";
            when "11" & x"efd" => data <= x"65";
            when "11" & x"efe" => data <= x"c4";
            when "11" & x"eff" => data <= x"85";
            when "11" & x"f00" => data <= x"c4";
            when "11" & x"f01" => data <= x"90";
            when "11" & x"f02" => data <= x"02";
            when "11" & x"f03" => data <= x"e6";
            when "11" & x"f04" => data <= x"c5";
            when "11" & x"f05" => data <= x"c8";
            when "11" & x"f06" => data <= x"b1";
            when "11" & x"f07" => data <= x"b0";
            when "11" & x"f08" => data <= x"c9";
            when "11" & x"f09" => data <= x"0a";
            when "11" & x"f0a" => data <= x"b0";
            when "11" & x"f0b" => data <= x"95";
            when "11" & x"f0c" => data <= x"18";
            when "11" & x"f0d" => data <= x"65";
            when "11" & x"f0e" => data <= x"c4";
            when "11" & x"f0f" => data <= x"85";
            when "11" & x"f10" => data <= x"c4";
            when "11" & x"f11" => data <= x"90";
            when "11" & x"f12" => data <= x"02";
            when "11" & x"f13" => data <= x"e6";
            when "11" & x"f14" => data <= x"c5";
            when "11" & x"f15" => data <= x"18";
            when "11" & x"f16" => data <= x"a9";
            when "11" & x"f17" => data <= x"00";
            when "11" & x"f18" => data <= x"8d";
            when "11" & x"f19" => data <= x"28";
            when "11" & x"f1a" => data <= x"0d";
            when "11" & x"f1b" => data <= x"a5";
            when "11" & x"f1c" => data <= x"c5";
            when "11" & x"f1d" => data <= x"6a";
            when "11" & x"f1e" => data <= x"48";
            when "11" & x"f1f" => data <= x"a5";
            when "11" & x"f20" => data <= x"c4";
            when "11" & x"f21" => data <= x"6a";
            when "11" & x"f22" => data <= x"48";
            when "11" & x"f23" => data <= x"90";
            when "11" & x"f24" => data <= x"03";
            when "11" & x"f25" => data <= x"6e";
            when "11" & x"f26" => data <= x"28";
            when "11" & x"f27" => data <= x"0d";
            when "11" & x"f28" => data <= x"c8";
            when "11" & x"f29" => data <= x"b1";
            when "11" & x"f2a" => data <= x"b0";
            when "11" & x"f2b" => data <= x"29";
            when "11" & x"f2c" => data <= x"1f";
            when "11" & x"f2d" => data <= x"8d";
            when "11" & x"f2e" => data <= x"27";
            when "11" & x"f2f" => data <= x"0d";
            when "11" & x"f30" => data <= x"f0";
            when "11" & x"f31" => data <= x"55";
            when "11" & x"f32" => data <= x"18";
            when "11" & x"f33" => data <= x"65";
            when "11" & x"f34" => data <= x"c4";
            when "11" & x"f35" => data <= x"aa";
            when "11" & x"f36" => data <= x"a9";
            when "11" & x"f37" => data <= x"00";
            when "11" & x"f38" => data <= x"65";
            when "11" & x"f39" => data <= x"c5";
            when "11" & x"f3a" => data <= x"c9";
            when "11" & x"f3b" => data <= x"03";
            when "11" & x"f3c" => data <= x"90";
            when "11" & x"f3d" => data <= x"06";
            when "11" & x"f3e" => data <= x"d0";
            when "11" & x"f3f" => data <= x"51";
            when "11" & x"f40" => data <= x"e0";
            when "11" & x"f41" => data <= x"21";
            when "11" & x"f42" => data <= x"b0";
            when "11" & x"f43" => data <= x"4d";
            when "11" & x"f44" => data <= x"a6";
            when "11" & x"f45" => data <= x"c0";
            when "11" & x"f46" => data <= x"bd";
            when "11" & x"f47" => data <= x"10";
            when "11" & x"f48" => data <= x"0d";
            when "11" & x"f49" => data <= x"6a";
            when "11" & x"f4a" => data <= x"bd";
            when "11" & x"f4b" => data <= x"0c";
            when "11" & x"f4c" => data <= x"0d";
            when "11" & x"f4d" => data <= x"20";
            when "11" & x"f4e" => data <= x"26";
            when "11" & x"f4f" => data <= x"ae";
            when "11" & x"f50" => data <= x"18";
            when "11" & x"f51" => data <= x"68";
            when "11" & x"f52" => data <= x"6d";
            when "11" & x"f53" => data <= x"23";
            when "11" & x"f54" => data <= x"0d";
            when "11" & x"f55" => data <= x"8d";
            when "11" & x"f56" => data <= x"23";
            when "11" & x"f57" => data <= x"0d";
            when "11" & x"f58" => data <= x"68";
            when "11" & x"f59" => data <= x"6d";
            when "11" & x"f5a" => data <= x"24";
            when "11" & x"f5b" => data <= x"0d";
            when "11" & x"f5c" => data <= x"8d";
            when "11" & x"f5d" => data <= x"24";
            when "11" & x"f5e" => data <= x"0d";
            when "11" & x"f5f" => data <= x"ad";
            when "11" & x"f60" => data <= x"25";
            when "11" & x"f61" => data <= x"0d";
            when "11" & x"f62" => data <= x"69";
            when "11" & x"f63" => data <= x"00";
            when "11" & x"f64" => data <= x"8d";
            when "11" & x"f65" => data <= x"25";
            when "11" & x"f66" => data <= x"0d";
            when "11" & x"f67" => data <= x"ad";
            when "11" & x"f68" => data <= x"26";
            when "11" & x"f69" => data <= x"0d";
            when "11" & x"f6a" => data <= x"69";
            when "11" & x"f6b" => data <= x"00";
            when "11" & x"f6c" => data <= x"8d";
            when "11" & x"f6d" => data <= x"26";
            when "11" & x"f6e" => data <= x"0d";
            when "11" & x"f6f" => data <= x"a0";
            when "11" & x"f70" => data <= x"00";
            when "11" & x"f71" => data <= x"8c";
            when "11" & x"f72" => data <= x"29";
            when "11" & x"f73" => data <= x"0d";
            when "11" & x"f74" => data <= x"c8";
            when "11" & x"f75" => data <= x"b1";
            when "11" & x"f76" => data <= x"b0";
            when "11" & x"f77" => data <= x"85";
            when "11" & x"f78" => data <= x"a0";
            when "11" & x"f79" => data <= x"c8";
            when "11" & x"f7a" => data <= x"b1";
            when "11" & x"f7b" => data <= x"b0";
            when "11" & x"f7c" => data <= x"85";
            when "11" & x"f7d" => data <= x"a1";
            when "11" & x"f7e" => data <= x"a5";
            when "11" & x"f7f" => data <= x"bf";
            when "11" & x"f80" => data <= x"c9";
            when "11" & x"f81" => data <= x"13";
            when "11" & x"f82" => data <= x"f0";
            when "11" & x"f83" => data <= x"05";
            when "11" & x"f84" => data <= x"20";
            when "11" & x"f85" => data <= x"9f";
            when "11" & x"f86" => data <= x"af";
            when "11" & x"f87" => data <= x"18";
            when "11" & x"f88" => data <= x"60";
            when "11" & x"f89" => data <= x"20";
            when "11" & x"f8a" => data <= x"cc";
            when "11" & x"f8b" => data <= x"a7";
            when "11" & x"f8c" => data <= x"20";
            when "11" & x"f8d" => data <= x"cd";
            when "11" & x"f8e" => data <= x"a0";
            when "11" & x"f8f" => data <= x"18";
            when "11" & x"f90" => data <= x"60";
            when "11" & x"f91" => data <= x"a9";
            when "11" & x"f92" => data <= x"1e";
            when "11" & x"f93" => data <= x"38";
            when "11" & x"f94" => data <= x"60";
            when "11" & x"f95" => data <= x"44";
            when "11" & x"f96" => data <= x"55";
            when "11" & x"f97" => data <= x"49";
            when "11" & x"f98" => data <= x"4b";
            when "11" & x"f99" => data <= x"20";
            when "11" & x"f9a" => data <= x"44";
            when "11" & x"f9b" => data <= x"55";
            when "11" & x"f9c" => data <= x"49";
            when "11" & x"f9d" => data <= x"4b";
            when "11" & x"f9e" => data <= x"20";
            when "11" & x"f9f" => data <= x"44";
            when "11" & x"fa0" => data <= x"55";
            when "11" & x"fa1" => data <= x"49";
            when "11" & x"fa2" => data <= x"4b";
            when "11" & x"fa3" => data <= x"20";
            when "11" & x"fa4" => data <= x"44";
            when "11" & x"fa5" => data <= x"55";
            when "11" & x"fa6" => data <= x"49";
            when "11" & x"fa7" => data <= x"4b";
            when "11" & x"fa8" => data <= x"20";
            when "11" & x"fa9" => data <= x"44";
            when "11" & x"faa" => data <= x"55";
            when "11" & x"fab" => data <= x"49";
            when "11" & x"fac" => data <= x"4b";
            when "11" & x"fad" => data <= x"20";
            when "11" & x"fae" => data <= x"44";
            when "11" & x"faf" => data <= x"55";
            when "11" & x"fb0" => data <= x"49";
            when "11" & x"fb1" => data <= x"4b";
            when "11" & x"fb2" => data <= x"20";
            when "11" & x"fb3" => data <= x"44";
            when "11" & x"fb4" => data <= x"55";
            when "11" & x"fb5" => data <= x"49";
            when "11" & x"fb6" => data <= x"4b";
            when "11" & x"fb7" => data <= x"20";
            when "11" & x"fb8" => data <= x"44";
            when "11" & x"fb9" => data <= x"55";
            when "11" & x"fba" => data <= x"49";
            when "11" & x"fbb" => data <= x"4b";
            when "11" & x"fbc" => data <= x"20";
            when "11" & x"fbd" => data <= x"44";
            when "11" & x"fbe" => data <= x"55";
            when "11" & x"fbf" => data <= x"49";
            when "11" & x"fc0" => data <= x"4b";
            when "11" & x"fc1" => data <= x"20";
            when "11" & x"fc2" => data <= x"44";
            when "11" & x"fc3" => data <= x"55";
            when "11" & x"fc4" => data <= x"49";
            when "11" & x"fc5" => data <= x"4b";
            when "11" & x"fc6" => data <= x"20";
            when "11" & x"fc7" => data <= x"44";
            when "11" & x"fc8" => data <= x"55";
            when "11" & x"fc9" => data <= x"49";
            when "11" & x"fca" => data <= x"4b";
            when "11" & x"fcb" => data <= x"20";
            when "11" & x"fcc" => data <= x"44";
            when "11" & x"fcd" => data <= x"55";
            when "11" & x"fce" => data <= x"49";
            when "11" & x"fcf" => data <= x"4b";
            when "11" & x"fd0" => data <= x"20";
            when "11" & x"fd1" => data <= x"44";
            when "11" & x"fd2" => data <= x"55";
            when "11" & x"fd3" => data <= x"49";
            when "11" & x"fd4" => data <= x"4b";
            when "11" & x"fd5" => data <= x"20";
            when "11" & x"fd6" => data <= x"44";
            when "11" & x"fd7" => data <= x"55";
            when "11" & x"fd8" => data <= x"49";
            when "11" & x"fd9" => data <= x"4b";
            when "11" & x"fda" => data <= x"20";
            when "11" & x"fdb" => data <= x"44";
            when "11" & x"fdc" => data <= x"55";
            when "11" & x"fdd" => data <= x"49";
            when "11" & x"fde" => data <= x"4b";
            when "11" & x"fdf" => data <= x"20";
            when "11" & x"fe0" => data <= x"44";
            when "11" & x"fe1" => data <= x"55";
            when "11" & x"fe2" => data <= x"49";
            when "11" & x"fe3" => data <= x"4b";
            when "11" & x"fe4" => data <= x"20";
            when "11" & x"fe5" => data <= x"44";
            when "11" & x"fe6" => data <= x"55";
            when "11" & x"fe7" => data <= x"49";
            when "11" & x"fe8" => data <= x"4b";
            when "11" & x"fe9" => data <= x"20";
            when "11" & x"fea" => data <= x"44";
            when "11" & x"feb" => data <= x"55";
            when "11" & x"fec" => data <= x"49";
            when "11" & x"fed" => data <= x"4b";
            when "11" & x"fee" => data <= x"20";
            when "11" & x"fef" => data <= x"44";
            when "11" & x"ff0" => data <= x"55";
            when "11" & x"ff1" => data <= x"49";
            when "11" & x"ff2" => data <= x"4b";
            when "11" & x"ff3" => data <= x"20";
            when "11" & x"ff4" => data <= x"44";
            when "11" & x"ff5" => data <= x"55";
            when "11" & x"ff6" => data <= x"49";
            when "11" & x"ff7" => data <= x"4b";
            when "11" & x"ff8" => data <= x"20";
            when "11" & x"ff9" => data <= x"44";
            when "11" & x"ffa" => data <= x"55";
            when "11" & x"ffb" => data <= x"49";
            when "11" & x"ffc" => data <= x"4b";
            when "11" & x"ffd" => data <= x"20";
            when "11" & x"ffe" => data <= x"44";
            when "11" & x"fff" => data <= x"00";
            when others => data <= (others => '0');
        end case;
    end process;
end RTL;
