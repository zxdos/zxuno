-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb9",
     9 => x"8c080b0b",
    10 => x"0bb99008",
    11 => x"0b0b0bb9",
    12 => x"94080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b9940c0b",
    16 => x"0b0bb990",
    17 => x"0c0b0b0b",
    18 => x"b98c0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb3b4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b98c7080",
    57 => x"c3c4278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188c904",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bb99c0c",
    65 => x"9f0bb9a0",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"b9a008ff",
    69 => x"05b9a00c",
    70 => x"b9a00880",
    71 => x"25eb38b9",
    72 => x"9c08ff05",
    73 => x"b99c0cb9",
    74 => x"9c088025",
    75 => x"d738800b",
    76 => x"b9a00c80",
    77 => x"0bb99c0c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bb99c08",
    97 => x"258f3882",
    98 => x"bd2db99c",
    99 => x"08ff05b9",
   100 => x"9c0c82ff",
   101 => x"04b99c08",
   102 => x"b9a00853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"b99c08a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134b9a0",
   111 => x"088105b9",
   112 => x"a00cb9a0",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bb9a00c",
   116 => x"b99c0881",
   117 => x"05b99c0c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134b9",
   122 => x"a0088105",
   123 => x"b9a00cb9",
   124 => x"a008a02e",
   125 => x"0981068e",
   126 => x"38800bb9",
   127 => x"a00cb99c",
   128 => x"088105b9",
   129 => x"9c0c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bb9a4",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bb9a40c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872b9",
   169 => x"a4088407",
   170 => x"b9a40c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb5f8",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"b9a40852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"b98c0c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d0402fc",
   217 => x"050dec51",
   218 => x"8a710c86",
   219 => x"b72d8271",
   220 => x"0c028405",
   221 => x"0d0402fc",
   222 => x"050dec51",
   223 => x"92710c86",
   224 => x"b72d8271",
   225 => x"0c028405",
   226 => x"0d04a00b",
   227 => x"ec0c86b7",
   228 => x"2d0480c0",
   229 => x"0bec0c86",
   230 => x"b72d0402",
   231 => x"dc050d80",
   232 => x"59878a2d",
   233 => x"810bec0c",
   234 => x"7a52b9a8",
   235 => x"51aad82d",
   236 => x"b98c0879",
   237 => x"2e80ee38",
   238 => x"b9ac0870",
   239 => x"f80c79ff",
   240 => x"12565955",
   241 => x"73792e8b",
   242 => x"38811874",
   243 => x"812a5558",
   244 => x"73f738f7",
   245 => x"18588159",
   246 => x"80752580",
   247 => x"c8387752",
   248 => x"7351848b",
   249 => x"2db9fc52",
   250 => x"b9a851ad",
   251 => x"972db98c",
   252 => x"08802e9a",
   253 => x"38b9fc57",
   254 => x"83fc5676",
   255 => x"70840558",
   256 => x"08e80cfc",
   257 => x"16567580",
   258 => x"25f13888",
   259 => x"9504b98c",
   260 => x"08598480",
   261 => x"55b9a851",
   262 => x"ace92dfc",
   263 => x"80158115",
   264 => x"555587d8",
   265 => x"04840bec",
   266 => x"0c78802e",
   267 => x"8d38b5fc",
   268 => x"518fc62d",
   269 => x"8dc92d88",
   270 => x"c004b6dc",
   271 => x"518fc62d",
   272 => x"78b98c0c",
   273 => x"02a4050d",
   274 => x"0402f005",
   275 => x"0d840bec",
   276 => x"0c8d972d",
   277 => x"89e62d81",
   278 => x"f82d8352",
   279 => x"8cfc2d81",
   280 => x"5184f02d",
   281 => x"ff125271",
   282 => x"8025f138",
   283 => x"840bec0c",
   284 => x"b4ac5185",
   285 => x"fe2da1d7",
   286 => x"2db98c08",
   287 => x"802e80d1",
   288 => x"38879b51",
   289 => x"b3ac2db5",
   290 => x"fc518fc6",
   291 => x"2d8db62d",
   292 => x"89f22d8f",
   293 => x"d62db690",
   294 => x"0b80f52d",
   295 => x"b7c80870",
   296 => x"81065455",
   297 => x"5371802e",
   298 => x"85387281",
   299 => x"07537381",
   300 => x"2a708106",
   301 => x"51527180",
   302 => x"2e853872",
   303 => x"82075372",
   304 => x"fc0c8652",
   305 => x"b98c0883",
   306 => x"38845271",
   307 => x"ec0c8990",
   308 => x"04800bb9",
   309 => x"8c0c0290",
   310 => x"050d0471",
   311 => x"980c04ff",
   312 => x"b008b98c",
   313 => x"0c04810b",
   314 => x"ffb00c04",
   315 => x"800bffb0",
   316 => x"0c0402f4",
   317 => x"050d8af4",
   318 => x"04b98c08",
   319 => x"81f02e09",
   320 => x"81068938",
   321 => x"810bb7c0",
   322 => x"0c8af404",
   323 => x"b98c0881",
   324 => x"e02e0981",
   325 => x"06893881",
   326 => x"0bb7c40c",
   327 => x"8af404b9",
   328 => x"8c0852b7",
   329 => x"c408802e",
   330 => x"8838b98c",
   331 => x"08818005",
   332 => x"5271842c",
   333 => x"728f0653",
   334 => x"53b7c008",
   335 => x"802e9938",
   336 => x"728429b7",
   337 => x"80057213",
   338 => x"81712b70",
   339 => x"09730806",
   340 => x"730c5153",
   341 => x"538aea04",
   342 => x"728429b7",
   343 => x"80057213",
   344 => x"83712b72",
   345 => x"0807720c",
   346 => x"5353800b",
   347 => x"b7c40c80",
   348 => x"0bb7c00c",
   349 => x"b9b4518b",
   350 => x"f52db98c",
   351 => x"08ff24fe",
   352 => x"f838800b",
   353 => x"b98c0c02",
   354 => x"8c050d04",
   355 => x"02f8050d",
   356 => x"b780528f",
   357 => x"51807270",
   358 => x"8405540c",
   359 => x"ff115170",
   360 => x"8025f238",
   361 => x"0288050d",
   362 => x"0402f005",
   363 => x"0d755189",
   364 => x"ec2d7082",
   365 => x"2cfc06b7",
   366 => x"80117210",
   367 => x"9e067108",
   368 => x"70722a70",
   369 => x"83068274",
   370 => x"2b700974",
   371 => x"06760c54",
   372 => x"51565753",
   373 => x"515389e6",
   374 => x"2d71b98c",
   375 => x"0c029005",
   376 => x"0d0402fc",
   377 => x"050d7251",
   378 => x"80710c80",
   379 => x"0b84120c",
   380 => x"0284050d",
   381 => x"0402f005",
   382 => x"0d757008",
   383 => x"84120853",
   384 => x"5353ff54",
   385 => x"71712ea8",
   386 => x"3889ec2d",
   387 => x"84130870",
   388 => x"84291488",
   389 => x"11700870",
   390 => x"81ff0684",
   391 => x"18088111",
   392 => x"8706841a",
   393 => x"0c535155",
   394 => x"51515189",
   395 => x"e62d7154",
   396 => x"73b98c0c",
   397 => x"0290050d",
   398 => x"0402f805",
   399 => x"0d89ec2d",
   400 => x"e008708b",
   401 => x"2a708106",
   402 => x"51525270",
   403 => x"802e9d38",
   404 => x"b9b40870",
   405 => x"8429b9bc",
   406 => x"057381ff",
   407 => x"06710c51",
   408 => x"51b9b408",
   409 => x"81118706",
   410 => x"b9b40c51",
   411 => x"800bb9dc",
   412 => x"0c89df2d",
   413 => x"89e62d02",
   414 => x"88050d04",
   415 => x"02fc050d",
   416 => x"89ec2d81",
   417 => x"0bb9dc0c",
   418 => x"89e62db9",
   419 => x"dc085170",
   420 => x"fa380284",
   421 => x"050d0402",
   422 => x"fc050db9",
   423 => x"b4518be2",
   424 => x"2d8b8c2d",
   425 => x"8cb95189",
   426 => x"db2d0284",
   427 => x"050d04b9",
   428 => x"e808b98c",
   429 => x"0c0402fc",
   430 => x"050d810b",
   431 => x"b7cc0c81",
   432 => x"5184f02d",
   433 => x"0284050d",
   434 => x"0402fc05",
   435 => x"0d8dd304",
   436 => x"89f22d80",
   437 => x"f6518ba9",
   438 => x"2db98c08",
   439 => x"f33880da",
   440 => x"518ba92d",
   441 => x"b98c08e8",
   442 => x"38b98c08",
   443 => x"b7cc0cb9",
   444 => x"8c085184",
   445 => x"f02d0284",
   446 => x"050d0402",
   447 => x"ec050d76",
   448 => x"54805287",
   449 => x"0b881580",
   450 => x"f52d5653",
   451 => x"74722483",
   452 => x"38a05372",
   453 => x"5182f92d",
   454 => x"81128b15",
   455 => x"80f52d54",
   456 => x"52727225",
   457 => x"de380294",
   458 => x"050d0402",
   459 => x"f0050db9",
   460 => x"e8085481",
   461 => x"f82d800b",
   462 => x"b9ec0c73",
   463 => x"08802e81",
   464 => x"8038820b",
   465 => x"b9a00cb9",
   466 => x"ec088f06",
   467 => x"b99c0c73",
   468 => x"08527183",
   469 => x"2e963871",
   470 => x"83268938",
   471 => x"71812eaf",
   472 => x"388fac04",
   473 => x"71852e9f",
   474 => x"388fac04",
   475 => x"881480f5",
   476 => x"2d841508",
   477 => x"b4c45354",
   478 => x"5285fe2d",
   479 => x"71842913",
   480 => x"70085252",
   481 => x"8fb00473",
   482 => x"518dfb2d",
   483 => x"8fac04b7",
   484 => x"c8088815",
   485 => x"082c7081",
   486 => x"06515271",
   487 => x"802e8738",
   488 => x"b4c8518f",
   489 => x"a904b4cc",
   490 => x"5185fe2d",
   491 => x"84140851",
   492 => x"85fe2db9",
   493 => x"ec088105",
   494 => x"b9ec0c8c",
   495 => x"14548ebb",
   496 => x"04029005",
   497 => x"0d0471b9",
   498 => x"e80c8eab",
   499 => x"2db9ec08",
   500 => x"ff05b9f0",
   501 => x"0c0402e8",
   502 => x"050db9e8",
   503 => x"08b9f408",
   504 => x"575580f6",
   505 => x"518ba92d",
   506 => x"b98c0881",
   507 => x"2a708106",
   508 => x"51527180",
   509 => x"2ea1388f",
   510 => x"fd0489f2",
   511 => x"2d80f651",
   512 => x"8ba92db9",
   513 => x"8c08f338",
   514 => x"b7cc0881",
   515 => x"3270b7cc",
   516 => x"0c705252",
   517 => x"84f02d80",
   518 => x"0bb9e00c",
   519 => x"800bb9e4",
   520 => x"0cb7cc08",
   521 => x"83b93880",
   522 => x"da518ba9",
   523 => x"2db98c08",
   524 => x"802e8a38",
   525 => x"b9e00881",
   526 => x"8007b9e0",
   527 => x"0c80d951",
   528 => x"8ba92db9",
   529 => x"8c08802e",
   530 => x"8a38b9e0",
   531 => x"0880c007",
   532 => x"b9e00c81",
   533 => x"94518ba9",
   534 => x"2db98c08",
   535 => x"802e8938",
   536 => x"b9e00890",
   537 => x"07b9e00c",
   538 => x"8191518b",
   539 => x"a92db98c",
   540 => x"08802e89",
   541 => x"38b9e008",
   542 => x"a007b9e0",
   543 => x"0c81f551",
   544 => x"8ba92db9",
   545 => x"8c08802e",
   546 => x"8938b9e0",
   547 => x"088107b9",
   548 => x"e00c81f2",
   549 => x"518ba92d",
   550 => x"b98c0880",
   551 => x"2e8938b9",
   552 => x"e0088207",
   553 => x"b9e00c81",
   554 => x"eb518ba9",
   555 => x"2db98c08",
   556 => x"802e8938",
   557 => x"b9e00884",
   558 => x"07b9e00c",
   559 => x"81f4518b",
   560 => x"a92db98c",
   561 => x"08802e89",
   562 => x"38b9e008",
   563 => x"8807b9e0",
   564 => x"0c80d851",
   565 => x"8ba92db9",
   566 => x"8c08802e",
   567 => x"8a38b9e4",
   568 => x"08818007",
   569 => x"b9e40c92",
   570 => x"518ba92d",
   571 => x"b98c0880",
   572 => x"2e8a38b9",
   573 => x"e40880c0",
   574 => x"07b9e40c",
   575 => x"94518ba9",
   576 => x"2db98c08",
   577 => x"802e8938",
   578 => x"b9e40890",
   579 => x"07b9e40c",
   580 => x"91518ba9",
   581 => x"2db98c08",
   582 => x"802e8938",
   583 => x"b9e408a0",
   584 => x"07b9e40c",
   585 => x"9d518ba9",
   586 => x"2db98c08",
   587 => x"802e8938",
   588 => x"b9e40881",
   589 => x"07b9e40c",
   590 => x"9b518ba9",
   591 => x"2db98c08",
   592 => x"802e8938",
   593 => x"b9e40882",
   594 => x"07b9e40c",
   595 => x"9c518ba9",
   596 => x"2db98c08",
   597 => x"802e8938",
   598 => x"b9e40884",
   599 => x"07b9e40c",
   600 => x"a3518ba9",
   601 => x"2db98c08",
   602 => x"802e8938",
   603 => x"b9e40888",
   604 => x"07b9e40c",
   605 => x"96518ba9",
   606 => x"2db98c08",
   607 => x"802e8438",
   608 => x"86f62d9e",
   609 => x"518ba92d",
   610 => x"b98c0880",
   611 => x"2e843886",
   612 => x"e22d9451",
   613 => x"8ba92db9",
   614 => x"8c088e38",
   615 => x"8194518b",
   616 => x"a92db98c",
   617 => x"08802ea8",
   618 => x"3891518b",
   619 => x"a92db98c",
   620 => x"088e3881",
   621 => x"91518ba9",
   622 => x"2db98c08",
   623 => x"802e9138",
   624 => x"80e6518b",
   625 => x"a92db98c",
   626 => x"08802e84",
   627 => x"3887922d",
   628 => x"81fd518b",
   629 => x"a92d81fa",
   630 => x"518ba92d",
   631 => x"99ce0494",
   632 => x"518ba92d",
   633 => x"b98c088e",
   634 => x"38819451",
   635 => x"8ba92db9",
   636 => x"8c08802e",
   637 => x"a8389151",
   638 => x"8ba92db9",
   639 => x"8c088e38",
   640 => x"8191518b",
   641 => x"a92db98c",
   642 => x"08802e91",
   643 => x"3880e651",
   644 => x"8ba92db9",
   645 => x"8c08802e",
   646 => x"84388792",
   647 => x"2d81f551",
   648 => x"8ba92db9",
   649 => x"8c08812a",
   650 => x"70810651",
   651 => x"5271802e",
   652 => x"af38b9f0",
   653 => x"08527180",
   654 => x"2e8938ff",
   655 => x"12b9f00c",
   656 => x"94e004b9",
   657 => x"ec0810b9",
   658 => x"ec080570",
   659 => x"84291651",
   660 => x"52881208",
   661 => x"802e8938",
   662 => x"ff518812",
   663 => x"0852712d",
   664 => x"81f2518b",
   665 => x"a92db98c",
   666 => x"08812a70",
   667 => x"81065152",
   668 => x"71802eb1",
   669 => x"38b9ec08",
   670 => x"ff11b9f0",
   671 => x"08565353",
   672 => x"73722589",
   673 => x"388114b9",
   674 => x"f00c95a5",
   675 => x"04721013",
   676 => x"70842916",
   677 => x"51528812",
   678 => x"08802e89",
   679 => x"38fe5188",
   680 => x"12085271",
   681 => x"2d81fd51",
   682 => x"8ba92db9",
   683 => x"8c08812a",
   684 => x"70810651",
   685 => x"5271802e",
   686 => x"ad38b9f0",
   687 => x"08802e89",
   688 => x"38800bb9",
   689 => x"f00c95e6",
   690 => x"04b9ec08",
   691 => x"10b9ec08",
   692 => x"05708429",
   693 => x"16515288",
   694 => x"1208802e",
   695 => x"8938fd51",
   696 => x"88120852",
   697 => x"712d81fa",
   698 => x"518ba92d",
   699 => x"b98c0881",
   700 => x"2a708106",
   701 => x"51527180",
   702 => x"2eae38b9",
   703 => x"ec08ff11",
   704 => x"5452b9f0",
   705 => x"08732588",
   706 => x"3872b9f0",
   707 => x"0c96a804",
   708 => x"71101270",
   709 => x"84291651",
   710 => x"52881208",
   711 => x"802e8938",
   712 => x"fc518812",
   713 => x"0852712d",
   714 => x"b9f00870",
   715 => x"53547380",
   716 => x"2e8a388c",
   717 => x"15ff1555",
   718 => x"5596ae04",
   719 => x"820bb9a0",
   720 => x"0c718f06",
   721 => x"b99c0c81",
   722 => x"eb518ba9",
   723 => x"2db98c08",
   724 => x"812a7081",
   725 => x"06515271",
   726 => x"802ead38",
   727 => x"7408852e",
   728 => x"098106a4",
   729 => x"38881580",
   730 => x"f52dff05",
   731 => x"52718816",
   732 => x"81b72d71",
   733 => x"982b5271",
   734 => x"80258838",
   735 => x"800b8816",
   736 => x"81b72d74",
   737 => x"518dfb2d",
   738 => x"81f4518b",
   739 => x"a92db98c",
   740 => x"08812a70",
   741 => x"81065152",
   742 => x"71802eb3",
   743 => x"38740885",
   744 => x"2e098106",
   745 => x"aa388815",
   746 => x"80f52d81",
   747 => x"05527188",
   748 => x"1681b72d",
   749 => x"7181ff06",
   750 => x"8b1680f5",
   751 => x"2d545272",
   752 => x"72278738",
   753 => x"72881681",
   754 => x"b72d7451",
   755 => x"8dfb2d80",
   756 => x"da518ba9",
   757 => x"2db98c08",
   758 => x"812a7081",
   759 => x"06515271",
   760 => x"802e81a6",
   761 => x"38b9e808",
   762 => x"b9f00855",
   763 => x"5373802e",
   764 => x"8a388c13",
   765 => x"ff155553",
   766 => x"97ed0472",
   767 => x"08527182",
   768 => x"2ea63871",
   769 => x"82268938",
   770 => x"71812ea9",
   771 => x"38998a04",
   772 => x"71832eb1",
   773 => x"3871842e",
   774 => x"09810680",
   775 => x"ed388813",
   776 => x"08518fc6",
   777 => x"2d998a04",
   778 => x"b9f00851",
   779 => x"88130852",
   780 => x"712d998a",
   781 => x"04810b88",
   782 => x"14082bb7",
   783 => x"c80832b7",
   784 => x"c80c98e0",
   785 => x"04881380",
   786 => x"f52d8105",
   787 => x"8b1480f5",
   788 => x"2d535471",
   789 => x"74248338",
   790 => x"80547388",
   791 => x"1481b72d",
   792 => x"8eab2d99",
   793 => x"8a047508",
   794 => x"802ea238",
   795 => x"7508518b",
   796 => x"a92db98c",
   797 => x"08810652",
   798 => x"71802e8b",
   799 => x"38b9f008",
   800 => x"51841608",
   801 => x"52712d88",
   802 => x"165675da",
   803 => x"38805480",
   804 => x"0bb9a00c",
   805 => x"738f06b9",
   806 => x"9c0ca052",
   807 => x"73b9f008",
   808 => x"2e098106",
   809 => x"9838b9ec",
   810 => x"08ff0574",
   811 => x"32700981",
   812 => x"05707207",
   813 => x"9f2a9171",
   814 => x"31515153",
   815 => x"53715182",
   816 => x"f92d8114",
   817 => x"548e7425",
   818 => x"c638b7cc",
   819 => x"085271b9",
   820 => x"8c0c0298",
   821 => x"050d0402",
   822 => x"f4050dd4",
   823 => x"5281ff72",
   824 => x"0c710853",
   825 => x"81ff720c",
   826 => x"72882b83",
   827 => x"fe800672",
   828 => x"087081ff",
   829 => x"06515253",
   830 => x"81ff720c",
   831 => x"72710788",
   832 => x"2b720870",
   833 => x"81ff0651",
   834 => x"525381ff",
   835 => x"720c7271",
   836 => x"07882b72",
   837 => x"087081ff",
   838 => x"067207b9",
   839 => x"8c0c5253",
   840 => x"028c050d",
   841 => x"0402f405",
   842 => x"0d747671",
   843 => x"81ff06d4",
   844 => x"0c5353b9",
   845 => x"f8088538",
   846 => x"71892b52",
   847 => x"71982ad4",
   848 => x"0c71902a",
   849 => x"7081ff06",
   850 => x"d40c5171",
   851 => x"882a7081",
   852 => x"ff06d40c",
   853 => x"517181ff",
   854 => x"06d40c72",
   855 => x"902a7081",
   856 => x"ff06d40c",
   857 => x"51d40870",
   858 => x"81ff0651",
   859 => x"5182b8bf",
   860 => x"527081ff",
   861 => x"2e098106",
   862 => x"943881ff",
   863 => x"0bd40cd4",
   864 => x"087081ff",
   865 => x"06ff1454",
   866 => x"515171e5",
   867 => x"3870b98c",
   868 => x"0c028c05",
   869 => x"0d0402fc",
   870 => x"050d81c7",
   871 => x"5181ff0b",
   872 => x"d40cff11",
   873 => x"51708025",
   874 => x"f4380284",
   875 => x"050d0402",
   876 => x"f4050d81",
   877 => x"ff0bd40c",
   878 => x"93538052",
   879 => x"87fc80c1",
   880 => x"519aa52d",
   881 => x"b98c088b",
   882 => x"3881ff0b",
   883 => x"d40c8153",
   884 => x"9bdc049b",
   885 => x"962dff13",
   886 => x"5372df38",
   887 => x"72b98c0c",
   888 => x"028c050d",
   889 => x"0402ec05",
   890 => x"0d810bb9",
   891 => x"f80c8454",
   892 => x"d008708f",
   893 => x"2a708106",
   894 => x"51515372",
   895 => x"f33872d0",
   896 => x"0c9b962d",
   897 => x"b4d05185",
   898 => x"fe2dd008",
   899 => x"708f2a70",
   900 => x"81065151",
   901 => x"5372f338",
   902 => x"810bd00c",
   903 => x"b1538052",
   904 => x"84d480c0",
   905 => x"519aa52d",
   906 => x"b98c0881",
   907 => x"2e933872",
   908 => x"822ebd38",
   909 => x"ff135372",
   910 => x"e538ff14",
   911 => x"5473ffb0",
   912 => x"389b962d",
   913 => x"83aa5284",
   914 => x"9c80c851",
   915 => x"9aa52db9",
   916 => x"8c08812e",
   917 => x"09810692",
   918 => x"3899d72d",
   919 => x"b98c0883",
   920 => x"ffff0653",
   921 => x"7283aa2e",
   922 => x"9d389baf",
   923 => x"2d9d8104",
   924 => x"b4dc5185",
   925 => x"fe2d8053",
   926 => x"9ecf04b4",
   927 => x"f45185fe",
   928 => x"2d80549e",
   929 => x"a10481ff",
   930 => x"0bd40cb1",
   931 => x"549b962d",
   932 => x"8fcf5380",
   933 => x"5287fc80",
   934 => x"f7519aa5",
   935 => x"2db98c08",
   936 => x"55b98c08",
   937 => x"812e0981",
   938 => x"069b3881",
   939 => x"ff0bd40c",
   940 => x"820a5284",
   941 => x"9c80e951",
   942 => x"9aa52db9",
   943 => x"8c08802e",
   944 => x"8d389b96",
   945 => x"2dff1353",
   946 => x"72c9389e",
   947 => x"940481ff",
   948 => x"0bd40cb9",
   949 => x"8c085287",
   950 => x"fc80fa51",
   951 => x"9aa52db9",
   952 => x"8c08b138",
   953 => x"81ff0bd4",
   954 => x"0cd40853",
   955 => x"81ff0bd4",
   956 => x"0c81ff0b",
   957 => x"d40c81ff",
   958 => x"0bd40c81",
   959 => x"ff0bd40c",
   960 => x"72862a70",
   961 => x"81067656",
   962 => x"51537295",
   963 => x"38b98c08",
   964 => x"549ea104",
   965 => x"73822efe",
   966 => x"e238ff14",
   967 => x"5473feed",
   968 => x"3873b9f8",
   969 => x"0c738b38",
   970 => x"815287fc",
   971 => x"80d0519a",
   972 => x"a52d81ff",
   973 => x"0bd40cd0",
   974 => x"08708f2a",
   975 => x"70810651",
   976 => x"515372f3",
   977 => x"3872d00c",
   978 => x"81ff0bd4",
   979 => x"0c815372",
   980 => x"b98c0c02",
   981 => x"94050d04",
   982 => x"02e8050d",
   983 => x"78558056",
   984 => x"81ff0bd4",
   985 => x"0cd00870",
   986 => x"8f2a7081",
   987 => x"06515153",
   988 => x"72f33882",
   989 => x"810bd00c",
   990 => x"81ff0bd4",
   991 => x"0c775287",
   992 => x"fc80d151",
   993 => x"9aa52d80",
   994 => x"dbc6df54",
   995 => x"b98c0880",
   996 => x"2e8a38b5",
   997 => x"945185fe",
   998 => x"2d9fef04",
   999 => x"81ff0bd4",
  1000 => x"0cd40870",
  1001 => x"81ff0651",
  1002 => x"537281fe",
  1003 => x"2e098106",
  1004 => x"9d3880ff",
  1005 => x"5399d72d",
  1006 => x"b98c0875",
  1007 => x"70840557",
  1008 => x"0cff1353",
  1009 => x"728025ed",
  1010 => x"3881569f",
  1011 => x"d404ff14",
  1012 => x"5473c938",
  1013 => x"81ff0bd4",
  1014 => x"0c81ff0b",
  1015 => x"d40cd008",
  1016 => x"708f2a70",
  1017 => x"81065151",
  1018 => x"5372f338",
  1019 => x"72d00c75",
  1020 => x"b98c0c02",
  1021 => x"98050d04",
  1022 => x"02e8050d",
  1023 => x"77797b58",
  1024 => x"55558053",
  1025 => x"727625a3",
  1026 => x"38747081",
  1027 => x"055680f5",
  1028 => x"2d747081",
  1029 => x"055680f5",
  1030 => x"2d525271",
  1031 => x"712e8638",
  1032 => x"8151a0ad",
  1033 => x"04811353",
  1034 => x"a0840480",
  1035 => x"5170b98c",
  1036 => x"0c029805",
  1037 => x"0d0402ec",
  1038 => x"050d7655",
  1039 => x"74802ebe",
  1040 => x"389a1580",
  1041 => x"e02d51ad",
  1042 => x"f02db98c",
  1043 => x"08b98c08",
  1044 => x"80c0ac0c",
  1045 => x"b98c0854",
  1046 => x"5480c088",
  1047 => x"08802e99",
  1048 => x"38941580",
  1049 => x"e02d51ad",
  1050 => x"f02db98c",
  1051 => x"08902b83",
  1052 => x"fff00a06",
  1053 => x"70750751",
  1054 => x"537280c0",
  1055 => x"ac0c80c0",
  1056 => x"ac085372",
  1057 => x"802e9d38",
  1058 => x"80c08008",
  1059 => x"fe147129",
  1060 => x"80c09408",
  1061 => x"0580c0b0",
  1062 => x"0c70842b",
  1063 => x"80c08c0c",
  1064 => x"54a1d204",
  1065 => x"80c09808",
  1066 => x"80c0ac0c",
  1067 => x"80c09c08",
  1068 => x"80c0b00c",
  1069 => x"80c08808",
  1070 => x"802e8b38",
  1071 => x"80c08008",
  1072 => x"842b53a1",
  1073 => x"cd0480c0",
  1074 => x"a008842b",
  1075 => x"537280c0",
  1076 => x"8c0c0294",
  1077 => x"050d0402",
  1078 => x"d8050d80",
  1079 => x"0b80c088",
  1080 => x"0c84549b",
  1081 => x"e52db98c",
  1082 => x"08802e95",
  1083 => x"38b9fc52",
  1084 => x"80519ed8",
  1085 => x"2db98c08",
  1086 => x"802e8638",
  1087 => x"fe54a289",
  1088 => x"04ff1454",
  1089 => x"738024db",
  1090 => x"38738c38",
  1091 => x"b5a45185",
  1092 => x"fe2d7355",
  1093 => x"a7ab0480",
  1094 => x"56810b80",
  1095 => x"c0b40c88",
  1096 => x"53b5b852",
  1097 => x"bab2519f",
  1098 => x"f82db98c",
  1099 => x"08762e09",
  1100 => x"81068838",
  1101 => x"b98c0880",
  1102 => x"c0b40c88",
  1103 => x"53b5c452",
  1104 => x"bace519f",
  1105 => x"f82db98c",
  1106 => x"088838b9",
  1107 => x"8c0880c0",
  1108 => x"b40c80c0",
  1109 => x"b408802e",
  1110 => x"80f638bd",
  1111 => x"c20b80f5",
  1112 => x"2dbdc30b",
  1113 => x"80f52d71",
  1114 => x"982b7190",
  1115 => x"2b07bdc4",
  1116 => x"0b80f52d",
  1117 => x"70882b72",
  1118 => x"07bdc50b",
  1119 => x"80f52d71",
  1120 => x"07bdfa0b",
  1121 => x"80f52dbd",
  1122 => x"fb0b80f5",
  1123 => x"2d71882b",
  1124 => x"07535f54",
  1125 => x"525a5657",
  1126 => x"557381ab",
  1127 => x"aa2e0981",
  1128 => x"068d3875",
  1129 => x"51adc02d",
  1130 => x"b98c0856",
  1131 => x"a3bc0473",
  1132 => x"82d4d52e",
  1133 => x"8738b5d0",
  1134 => x"51a3fe04",
  1135 => x"b9fc5275",
  1136 => x"519ed82d",
  1137 => x"b98c0855",
  1138 => x"b98c0880",
  1139 => x"2e83dc38",
  1140 => x"8853b5c4",
  1141 => x"52bace51",
  1142 => x"9ff82db9",
  1143 => x"8c088a38",
  1144 => x"810b80c0",
  1145 => x"880ca484",
  1146 => x"048853b5",
  1147 => x"b852bab2",
  1148 => x"519ff82d",
  1149 => x"b98c0880",
  1150 => x"2e8a38b5",
  1151 => x"e45185fe",
  1152 => x"2da4de04",
  1153 => x"bdfa0b80",
  1154 => x"f52d5473",
  1155 => x"80d52e09",
  1156 => x"810680ca",
  1157 => x"38bdfb0b",
  1158 => x"80f52d54",
  1159 => x"7381aa2e",
  1160 => x"098106ba",
  1161 => x"38800bb9",
  1162 => x"fc0b80f5",
  1163 => x"2d565474",
  1164 => x"81e92e83",
  1165 => x"38815474",
  1166 => x"81eb2e8c",
  1167 => x"38805573",
  1168 => x"752e0981",
  1169 => x"0682e438",
  1170 => x"ba870b80",
  1171 => x"f52d5574",
  1172 => x"8d38ba88",
  1173 => x"0b80f52d",
  1174 => x"5473822e",
  1175 => x"86388055",
  1176 => x"a7ab04ba",
  1177 => x"890b80f5",
  1178 => x"2d7080c0",
  1179 => x"800cff05",
  1180 => x"80c0840c",
  1181 => x"ba8a0b80",
  1182 => x"f52dba8b",
  1183 => x"0b80f52d",
  1184 => x"58760577",
  1185 => x"82802905",
  1186 => x"7080c090",
  1187 => x"0cba8c0b",
  1188 => x"80f52d70",
  1189 => x"80c0a40c",
  1190 => x"80c08808",
  1191 => x"59575876",
  1192 => x"802e81ac",
  1193 => x"388853b5",
  1194 => x"c452bace",
  1195 => x"519ff82d",
  1196 => x"b98c0881",
  1197 => x"f63880c0",
  1198 => x"80087084",
  1199 => x"2b80c08c",
  1200 => x"0c7080c0",
  1201 => x"a00cbaa1",
  1202 => x"0b80f52d",
  1203 => x"baa00b80",
  1204 => x"f52d7182",
  1205 => x"802905ba",
  1206 => x"a20b80f5",
  1207 => x"2d708480",
  1208 => x"802912ba",
  1209 => x"a30b80f5",
  1210 => x"2d708180",
  1211 => x"0a291270",
  1212 => x"80c0a80c",
  1213 => x"80c0a408",
  1214 => x"712980c0",
  1215 => x"90080570",
  1216 => x"80c0940c",
  1217 => x"baa90b80",
  1218 => x"f52dbaa8",
  1219 => x"0b80f52d",
  1220 => x"71828029",
  1221 => x"05baaa0b",
  1222 => x"80f52d70",
  1223 => x"84808029",
  1224 => x"12baab0b",
  1225 => x"80f52d70",
  1226 => x"982b81f0",
  1227 => x"0a067205",
  1228 => x"7080c098",
  1229 => x"0cfe117e",
  1230 => x"29770580",
  1231 => x"c09c0c52",
  1232 => x"59524354",
  1233 => x"5e515259",
  1234 => x"525d5759",
  1235 => x"57a7a404",
  1236 => x"ba8e0b80",
  1237 => x"f52dba8d",
  1238 => x"0b80f52d",
  1239 => x"71828029",
  1240 => x"057080c0",
  1241 => x"8c0c70a0",
  1242 => x"2983ff05",
  1243 => x"70892a70",
  1244 => x"80c0a00c",
  1245 => x"ba930b80",
  1246 => x"f52dba92",
  1247 => x"0b80f52d",
  1248 => x"71828029",
  1249 => x"057080c0",
  1250 => x"a80c7b71",
  1251 => x"291e7080",
  1252 => x"c09c0c7d",
  1253 => x"80c0980c",
  1254 => x"730580c0",
  1255 => x"940c555e",
  1256 => x"51515555",
  1257 => x"8051a0b6",
  1258 => x"2d815574",
  1259 => x"b98c0c02",
  1260 => x"a8050d04",
  1261 => x"02ec050d",
  1262 => x"7670872c",
  1263 => x"7180ff06",
  1264 => x"55565480",
  1265 => x"c088088a",
  1266 => x"3873882c",
  1267 => x"7481ff06",
  1268 => x"5455b9fc",
  1269 => x"5280c090",
  1270 => x"0815519e",
  1271 => x"d82db98c",
  1272 => x"0854b98c",
  1273 => x"08802eb4",
  1274 => x"3880c088",
  1275 => x"08802e98",
  1276 => x"38728429",
  1277 => x"b9fc0570",
  1278 => x"085253ad",
  1279 => x"c02db98c",
  1280 => x"08f00a06",
  1281 => x"53a89a04",
  1282 => x"7210b9fc",
  1283 => x"057080e0",
  1284 => x"2d5253ad",
  1285 => x"f02db98c",
  1286 => x"08537254",
  1287 => x"73b98c0c",
  1288 => x"0294050d",
  1289 => x"0402e005",
  1290 => x"0d797084",
  1291 => x"2c80c0b0",
  1292 => x"0805718f",
  1293 => x"06525553",
  1294 => x"728938b9",
  1295 => x"fc527351",
  1296 => x"9ed82d72",
  1297 => x"a029b9fc",
  1298 => x"05548074",
  1299 => x"80f52d56",
  1300 => x"5374732e",
  1301 => x"83388153",
  1302 => x"7481e52e",
  1303 => x"81ef3881",
  1304 => x"70740654",
  1305 => x"5872802e",
  1306 => x"81e3388b",
  1307 => x"1480f52d",
  1308 => x"70832a79",
  1309 => x"06585676",
  1310 => x"9838b7d0",
  1311 => x"08537288",
  1312 => x"3872bdfc",
  1313 => x"0b81b72d",
  1314 => x"76b7d00c",
  1315 => x"7353aacf",
  1316 => x"04758f2e",
  1317 => x"09810681",
  1318 => x"b438749f",
  1319 => x"068d29bd",
  1320 => x"ef115153",
  1321 => x"811480f5",
  1322 => x"2d737081",
  1323 => x"055581b7",
  1324 => x"2d831480",
  1325 => x"f52d7370",
  1326 => x"81055581",
  1327 => x"b72d8514",
  1328 => x"80f52d73",
  1329 => x"70810555",
  1330 => x"81b72d87",
  1331 => x"1480f52d",
  1332 => x"73708105",
  1333 => x"5581b72d",
  1334 => x"891480f5",
  1335 => x"2d737081",
  1336 => x"055581b7",
  1337 => x"2d8e1480",
  1338 => x"f52d7370",
  1339 => x"81055581",
  1340 => x"b72d9014",
  1341 => x"80f52d73",
  1342 => x"70810555",
  1343 => x"81b72d92",
  1344 => x"1480f52d",
  1345 => x"73708105",
  1346 => x"5581b72d",
  1347 => x"941480f5",
  1348 => x"2d737081",
  1349 => x"055581b7",
  1350 => x"2d961480",
  1351 => x"f52d7370",
  1352 => x"81055581",
  1353 => x"b72d9814",
  1354 => x"80f52d73",
  1355 => x"70810555",
  1356 => x"81b72d9c",
  1357 => x"1480f52d",
  1358 => x"73708105",
  1359 => x"5581b72d",
  1360 => x"9e1480f5",
  1361 => x"2d7381b7",
  1362 => x"2d77b7d0",
  1363 => x"0c805372",
  1364 => x"b98c0c02",
  1365 => x"a0050d04",
  1366 => x"02cc050d",
  1367 => x"7e605e5a",
  1368 => x"800b80c0",
  1369 => x"ac0880c0",
  1370 => x"b008595c",
  1371 => x"56805880",
  1372 => x"c08c0878",
  1373 => x"2e81b038",
  1374 => x"778f06a0",
  1375 => x"17575473",
  1376 => x"8f38b9fc",
  1377 => x"52765181",
  1378 => x"17579ed8",
  1379 => x"2db9fc56",
  1380 => x"807680f5",
  1381 => x"2d565474",
  1382 => x"742e8338",
  1383 => x"81547481",
  1384 => x"e52e80f7",
  1385 => x"38817075",
  1386 => x"06555c73",
  1387 => x"802e80eb",
  1388 => x"388b1680",
  1389 => x"f52d9806",
  1390 => x"597880df",
  1391 => x"388b537c",
  1392 => x"5275519f",
  1393 => x"f82db98c",
  1394 => x"0880d038",
  1395 => x"9c160851",
  1396 => x"adc02db9",
  1397 => x"8c08841b",
  1398 => x"0c9a1680",
  1399 => x"e02d51ad",
  1400 => x"f02db98c",
  1401 => x"08b98c08",
  1402 => x"881c0cb9",
  1403 => x"8c085555",
  1404 => x"80c08808",
  1405 => x"802e9838",
  1406 => x"941680e0",
  1407 => x"2d51adf0",
  1408 => x"2db98c08",
  1409 => x"902b83ff",
  1410 => x"f00a0670",
  1411 => x"16515473",
  1412 => x"881b0c78",
  1413 => x"7a0c7b54",
  1414 => x"ace00481",
  1415 => x"185880c0",
  1416 => x"8c087826",
  1417 => x"fed23880",
  1418 => x"c0880880",
  1419 => x"2eb0387a",
  1420 => x"51a7b42d",
  1421 => x"b98c08b9",
  1422 => x"8c0880ff",
  1423 => x"fffff806",
  1424 => x"555b7380",
  1425 => x"fffffff8",
  1426 => x"2e9438b9",
  1427 => x"8c08fe05",
  1428 => x"80c08008",
  1429 => x"2980c094",
  1430 => x"080557aa",
  1431 => x"ed048054",
  1432 => x"73b98c0c",
  1433 => x"02b4050d",
  1434 => x"0402f405",
  1435 => x"0d747008",
  1436 => x"8105710c",
  1437 => x"700880c0",
  1438 => x"84080653",
  1439 => x"53718e38",
  1440 => x"88130851",
  1441 => x"a7b42db9",
  1442 => x"8c088814",
  1443 => x"0c810bb9",
  1444 => x"8c0c028c",
  1445 => x"050d0402",
  1446 => x"f0050d75",
  1447 => x"881108fe",
  1448 => x"0580c080",
  1449 => x"082980c0",
  1450 => x"94081172",
  1451 => x"0880c084",
  1452 => x"08060579",
  1453 => x"55535454",
  1454 => x"9ed82d02",
  1455 => x"90050d04",
  1456 => x"02f4050d",
  1457 => x"7470882a",
  1458 => x"83fe8006",
  1459 => x"7072982a",
  1460 => x"0772882b",
  1461 => x"87fc8080",
  1462 => x"0673982b",
  1463 => x"81f00a06",
  1464 => x"71730707",
  1465 => x"b98c0c56",
  1466 => x"51535102",
  1467 => x"8c050d04",
  1468 => x"02f8050d",
  1469 => x"028e0580",
  1470 => x"f52d7488",
  1471 => x"2b077083",
  1472 => x"ffff06b9",
  1473 => x"8c0c5102",
  1474 => x"88050d04",
  1475 => x"02f4050d",
  1476 => x"74767853",
  1477 => x"54528071",
  1478 => x"25973872",
  1479 => x"70810554",
  1480 => x"80f52d72",
  1481 => x"70810554",
  1482 => x"81b72dff",
  1483 => x"115170eb",
  1484 => x"38807281",
  1485 => x"b72d028c",
  1486 => x"050d0402",
  1487 => x"e8050d77",
  1488 => x"56807056",
  1489 => x"54737624",
  1490 => x"b33880c0",
  1491 => x"8c08742e",
  1492 => x"ab387351",
  1493 => x"a8a52db9",
  1494 => x"8c08b98c",
  1495 => x"08098105",
  1496 => x"70b98c08",
  1497 => x"079f2a77",
  1498 => x"05811757",
  1499 => x"57535374",
  1500 => x"76248938",
  1501 => x"80c08c08",
  1502 => x"7426d738",
  1503 => x"72b98c0c",
  1504 => x"0298050d",
  1505 => x"0402f005",
  1506 => x"0db98808",
  1507 => x"1651aebb",
  1508 => x"2db98c08",
  1509 => x"802e9c38",
  1510 => x"8b53b98c",
  1511 => x"0852bdfc",
  1512 => x"51ae8c2d",
  1513 => x"80c0b808",
  1514 => x"5473802e",
  1515 => x"8638bdfc",
  1516 => x"51732d02",
  1517 => x"90050d04",
  1518 => x"02dc050d",
  1519 => x"80705a55",
  1520 => x"74b98808",
  1521 => x"25b13880",
  1522 => x"c08c0875",
  1523 => x"2ea93878",
  1524 => x"51a8a52d",
  1525 => x"b98c0809",
  1526 => x"810570b9",
  1527 => x"8c08079f",
  1528 => x"2a760581",
  1529 => x"1b5b5654",
  1530 => x"74b98808",
  1531 => x"25893880",
  1532 => x"c08c0879",
  1533 => x"26d93880",
  1534 => x"557880c0",
  1535 => x"8c082781",
  1536 => x"d1387851",
  1537 => x"a8a52db9",
  1538 => x"8c08802e",
  1539 => x"81a538b9",
  1540 => x"8c088b05",
  1541 => x"80f52d70",
  1542 => x"842a7081",
  1543 => x"06771078",
  1544 => x"842bbdfc",
  1545 => x"0b80f52d",
  1546 => x"5c5c5351",
  1547 => x"55567380",
  1548 => x"2e80c838",
  1549 => x"7416822b",
  1550 => x"b1f60bb7",
  1551 => x"dc120c54",
  1552 => x"77753110",
  1553 => x"80c0bc11",
  1554 => x"55569074",
  1555 => x"70810556",
  1556 => x"81b72da0",
  1557 => x"7481b72d",
  1558 => x"7681ff06",
  1559 => x"81165854",
  1560 => x"73802e89",
  1561 => x"389c53bd",
  1562 => x"fc52b0f3",
  1563 => x"048b53b9",
  1564 => x"8c085280",
  1565 => x"c0be1651",
  1566 => x"b1ab0474",
  1567 => x"16822baf",
  1568 => x"850bb7dc",
  1569 => x"120c5476",
  1570 => x"81ff0681",
  1571 => x"16585473",
  1572 => x"802e8938",
  1573 => x"9c53bdfc",
  1574 => x"52b1a204",
  1575 => x"8b53b98c",
  1576 => x"08527775",
  1577 => x"311080c0",
  1578 => x"bc055176",
  1579 => x"55ae8c2d",
  1580 => x"b1c70474",
  1581 => x"90297531",
  1582 => x"701080c0",
  1583 => x"bc055154",
  1584 => x"b98c0874",
  1585 => x"81b72d81",
  1586 => x"1959748b",
  1587 => x"24a338af",
  1588 => x"f9047490",
  1589 => x"29753170",
  1590 => x"1080c0bc",
  1591 => x"058c7731",
  1592 => x"57515480",
  1593 => x"7481b72d",
  1594 => x"9e14ff16",
  1595 => x"565474f3",
  1596 => x"3802a405",
  1597 => x"0d0402fc",
  1598 => x"050db988",
  1599 => x"081351ae",
  1600 => x"bb2db98c",
  1601 => x"08802e88",
  1602 => x"38b98c08",
  1603 => x"51a0b62d",
  1604 => x"800bb988",
  1605 => x"0cafb82d",
  1606 => x"8eab2d02",
  1607 => x"84050d04",
  1608 => x"02fc050d",
  1609 => x"725170fd",
  1610 => x"2ead3870",
  1611 => x"fd248a38",
  1612 => x"70fc2e80",
  1613 => x"c438b381",
  1614 => x"0470fe2e",
  1615 => x"b13870ff",
  1616 => x"2e098106",
  1617 => x"bc38b988",
  1618 => x"08517080",
  1619 => x"2eb338ff",
  1620 => x"11b9880c",
  1621 => x"b38104b9",
  1622 => x"8808f005",
  1623 => x"70b9880c",
  1624 => x"51708025",
  1625 => x"9c38800b",
  1626 => x"b9880cb3",
  1627 => x"8104b988",
  1628 => x"088105b9",
  1629 => x"880cb381",
  1630 => x"04b98808",
  1631 => x"9005b988",
  1632 => x"0cafb82d",
  1633 => x"8eab2d02",
  1634 => x"84050d04",
  1635 => x"02fc050d",
  1636 => x"800bb988",
  1637 => x"0cafb82d",
  1638 => x"8daf2db9",
  1639 => x"8c08b8f8",
  1640 => x"0cb7d451",
  1641 => x"8fc62d02",
  1642 => x"84050d04",
  1643 => x"7180c0b8",
  1644 => x"0c040000",
  1645 => x"00ffffff",
  1646 => x"ff00ffff",
  1647 => x"ffff00ff",
  1648 => x"ffffff00",
  1649 => x"52657365",
  1650 => x"74204e45",
  1651 => x"53000000",
  1652 => x"5363616e",
  1653 => x"6c696e65",
  1654 => x"73000000",
  1655 => x"48513258",
  1656 => x"2046696c",
  1657 => x"74657200",
  1658 => x"50312053",
  1659 => x"656c6563",
  1660 => x"74000000",
  1661 => x"50312053",
  1662 => x"74617274",
  1663 => x"00000000",
  1664 => x"4c6f6164",
  1665 => x"20524f4d",
  1666 => x"20100000",
  1667 => x"45786974",
  1668 => x"00000000",
  1669 => x"524f4d20",
  1670 => x"6c6f6164",
  1671 => x"696e6720",
  1672 => x"6661696c",
  1673 => x"65640000",
  1674 => x"4f4b0000",
  1675 => x"496e6974",
  1676 => x"69616c69",
  1677 => x"7a696e67",
  1678 => x"20534420",
  1679 => x"63617264",
  1680 => x"0a000000",
  1681 => x"16200000",
  1682 => x"14200000",
  1683 => x"15200000",
  1684 => x"53442069",
  1685 => x"6e69742e",
  1686 => x"2e2e0a00",
  1687 => x"53442063",
  1688 => x"61726420",
  1689 => x"72657365",
  1690 => x"74206661",
  1691 => x"696c6564",
  1692 => x"210a0000",
  1693 => x"53444843",
  1694 => x"20657272",
  1695 => x"6f72210a",
  1696 => x"00000000",
  1697 => x"57726974",
  1698 => x"65206661",
  1699 => x"696c6564",
  1700 => x"0a000000",
  1701 => x"52656164",
  1702 => x"20666169",
  1703 => x"6c65640a",
  1704 => x"00000000",
  1705 => x"43617264",
  1706 => x"20696e69",
  1707 => x"74206661",
  1708 => x"696c6564",
  1709 => x"0a000000",
  1710 => x"46415431",
  1711 => x"36202020",
  1712 => x"00000000",
  1713 => x"46415433",
  1714 => x"32202020",
  1715 => x"00000000",
  1716 => x"4e6f2070",
  1717 => x"61727469",
  1718 => x"74696f6e",
  1719 => x"20736967",
  1720 => x"0a000000",
  1721 => x"42616420",
  1722 => x"70617274",
  1723 => x"0a000000",
  1724 => x"4261636b",
  1725 => x"00000000",
  1726 => x"00000002",
  1727 => x"00000002",
  1728 => x"000019c4",
  1729 => x"0000034e",
  1730 => x"00000001",
  1731 => x"000019d0",
  1732 => x"00000000",
  1733 => x"00000001",
  1734 => x"000019dc",
  1735 => x"00000001",
  1736 => x"00000002",
  1737 => x"000019e8",
  1738 => x"00000362",
  1739 => x"00000002",
  1740 => x"000019f4",
  1741 => x"00000376",
  1742 => x"00000002",
  1743 => x"00001a00",
  1744 => x"0000198c",
  1745 => x"00000002",
  1746 => x"00001a0c",
  1747 => x"000006c9",
  1748 => x"00000000",
  1749 => x"00000000",
  1750 => x"00000000",
  1751 => x"00000004",
  1752 => x"00001a14",
  1753 => x"00001b5c",
  1754 => x"00000004",
  1755 => x"00001a28",
  1756 => x"00001afc",
  1757 => x"00000000",
  1758 => x"00000000",
  1759 => x"00000000",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000002",
  1782 => x"0000203c",
  1783 => x"00001785",
  1784 => x"00000002",
  1785 => x"0000205a",
  1786 => x"00001785",
  1787 => x"00000002",
  1788 => x"00002078",
  1789 => x"00001785",
  1790 => x"00000002",
  1791 => x"00002096",
  1792 => x"00001785",
  1793 => x"00000002",
  1794 => x"000020b4",
  1795 => x"00001785",
  1796 => x"00000002",
  1797 => x"000020d2",
  1798 => x"00001785",
  1799 => x"00000002",
  1800 => x"000020f0",
  1801 => x"00001785",
  1802 => x"00000002",
  1803 => x"0000210e",
  1804 => x"00001785",
  1805 => x"00000002",
  1806 => x"0000212c",
  1807 => x"00001785",
  1808 => x"00000002",
  1809 => x"0000214a",
  1810 => x"00001785",
  1811 => x"00000002",
  1812 => x"00002168",
  1813 => x"00001785",
  1814 => x"00000002",
  1815 => x"00002186",
  1816 => x"00001785",
  1817 => x"00000002",
  1818 => x"000021a4",
  1819 => x"00001785",
  1820 => x"00000004",
  1821 => x"00001af0",
  1822 => x"00000000",
  1823 => x"00000000",
  1824 => x"00000000",
  1825 => x"00001920",
  1826 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

