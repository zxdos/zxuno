-------------------------------------------------------------------------------
-- $Id: dac-c.vhd,v 1.1 2005/10/25 21:09:58 arnim Exp $
-------------------------------------------------------------------------------

configuration dac_rtl_c0 of dac is

  for rtl
  end for;

end dac_rtl_c0;
