-------------------------------------------------------------------------------
--
-- FPGA Colecovision
--
-- $Id: cv_por-c.vhd,v 1.3 2006/01/05 22:25:25 arnim Exp $
--
-------------------------------------------------------------------------------

configuration cv_por_rtl_c0 of cv_por is

  for cyclone
  end for;

end cv_por_rtl_c0;
