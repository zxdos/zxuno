-------------------------------------------------------------------------------
--
-- FPGA Colecovision
--
-- $Id: generic_ram.vhd,v 1.2 2006/01/05 23:31:32 arnim Exp $
--
-- Generic RTL flavour.
--
-- Characteristics of the synchronous RAM:
--   - memory is updated with rising clock edge
--   - no read-through-write capability
--
-------------------------------------------------------------------------------
--
-- Copyright (c) 2006, Arnim Laeuger (arnim.laeuger@gmx.net)
--
-- All rights reserved
--
-- Redistribution and use in source and synthezised forms, with or without
-- modification, are permitted provided that the following conditions are met:
--
-- Redistributions of source code must retain the above copyright notice,
-- this list of conditions and the following disclaimer.
--
-- Redistributions in synthesized form must reproduce the above copyright
-- notice, this list of conditions and the following disclaimer in the
-- documentation and/or other materials provided with the distribution.
--
-- Neither the name of the author nor the names of other contributors may
-- be used to endorse or promote products derived from this software without
-- specific prior written permission.
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
-- PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE
-- LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
-- CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
-- SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
-- INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
-- CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.
--
-- Please report bugs to the author, but before you do so, please
-- make sure that this is not a derivative work and that
-- you have the latest version of this file.
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity ram_init is

  generic (
    addr_width_g : integer := 10;
    data_width_g : integer := 8
  );
  port (
    clk_i : in  std_logic;
    a_i   : in  std_logic_vector(addr_width_g-1 downto 0);
    we_i  : in  std_logic;
    d_i   : in  std_logic_vector(data_width_g-1 downto 0);
    d_o   : out std_logic_vector(data_width_g-1 downto 0)
  );

end ram_init;


library ieee;
use ieee.numeric_std.all;

architecture rtl of ram_init is

  type mem_t is array (natural range 0 to 2**addr_width_g-1) of
    std_logic_vector(d_i'range);
  signal mem_q : mem_t := (
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0000
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0008
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0010
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0018
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0020
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0028
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0030
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0038
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0040
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0048
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0050
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0058
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0060
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0068
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0070
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0078
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0080
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0088
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0090
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0098
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0100
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0108
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0110
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0118
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0120
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0128
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0130
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0138
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0140
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0148
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0150
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0158
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0160
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0168
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0170
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0178
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0180
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0188
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0190
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0198
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0200
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0208
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0210
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0218
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0220
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0228
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0230
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0238
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0240
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0248
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0250
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0258
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0260
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0268
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0270
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0278
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0280
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0288
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0290
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0298
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0300
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0308
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0310
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0318
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0320
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0328
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0330
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0338
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0340
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0348
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0350
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0358
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0360
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0368
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0370
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0378
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0380
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0388
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0390
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0398
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0400
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0408
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0410
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0418
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0420
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0428
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0430
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0438
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0440
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0448
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0450
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0458
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0460
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0468
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0470
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0478
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0480
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0488
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0490
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0498
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0500
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0508
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0510
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0518
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0520
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0528
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0530
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0538
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0540
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0548
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0550
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0558
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0560
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0568
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0570
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0578
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0580
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0588
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0590
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0598
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05F8
    x"CD",x"E9",x"18",x"CD",x"85",x"1F",x"CD",x"D6", -- 0x0600
    x"1F",x"CD",x"97",x"77",x"21",x"00",x"20",x"3E", -- 0x0608
    x"F4",x"11",x"20",x"00",x"CD",x"82",x"1F",x"CD", -- 0x0610
    x"7F",x"1F",x"11",x"61",x"18",x"21",x"A6",x"77", -- 0x0618
    x"01",x"1C",x"00",x"CD",x"DF",x"1F",x"11",x"E1", -- 0x0620
    x"18",x"21",x"C2",x"77",x"01",x"1C",x"00",x"CD", -- 0x0628
    x"DF",x"1F",x"01",x"C2",x"01",x"CD",x"D9",x"1F", -- 0x0630
    x"21",x"01",x"00",x"CD",x"79",x"1F",x"7D",x"FE", -- 0x0638
    x"0F",x"28",x"F5",x"FE",x"0A",x"CA",x"4D",x"76", -- 0x0640
    x"FE",x"0B",x"C2",x"6E",x"00",x"11",x"E1",x"18", -- 0x0648
    x"21",x"DE",x"77",x"01",x"1C",x"00",x"CD",x"DF", -- 0x0650
    x"1F",x"3E",x"00",x"D3",x"21",x"3E",x"80",x"D3", -- 0x0658
    x"23",x"3E",x"23",x"D3",x"20",x"3E",x"00",x"D3", -- 0x0660
    x"21",x"3E",x"03",x"D3",x"23",x"3E",x"0B",x"D3", -- 0x0668
    x"24",x"C3",x"74",x"76",x"21",x"00",x"80",x"22", -- 0x0670
    x"A4",x"77",x"3E",x"00",x"32",x"A2",x"77",x"CD", -- 0x0678
    x"9C",x"76",x"DA",x"91",x"76",x"CD",x"57",x"77", -- 0x0680
    x"CD",x"4F",x"77",x"CD",x"2C",x"77",x"C3",x"7F", -- 0x0688
    x"76",x"CD",x"2C",x"77",x"3E",x"47",x"CD",x"8B", -- 0x0690
    x"77",x"C3",x"6E",x"00",x"AF",x"32",x"A3",x"77", -- 0x0698
    x"06",x"0A",x"CD",x"68",x"77",x"DA",x"D6",x"76", -- 0x06A0
    x"FE",x"01",x"CA",x"D9",x"76",x"B7",x"CA",x"A0", -- 0x06A8
    x"76",x"FE",x"04",x"37",x"C8",x"06",x"01",x"CD", -- 0x06B0
    x"68",x"77",x"D2",x"B5",x"76",x"3E",x"15",x"CD", -- 0x06B8
    x"8B",x"77",x"3A",x"A3",x"77",x"3C",x"32",x"A3", -- 0x06C0
    x"77",x"FE",x"0A",x"DA",x"A0",x"76",x"3E",x"45", -- 0x06C8
    x"CD",x"8B",x"77",x"C3",x"00",x"00",x"C3",x"B5", -- 0x06D0
    x"76",x"06",x"01",x"CD",x"68",x"77",x"DA",x"D6", -- 0x06D8
    x"76",x"57",x"06",x"01",x"CD",x"68",x"77",x"DA", -- 0x06E0
    x"D6",x"76",x"2F",x"BA",x"CA",x"F2",x"76",x"C3", -- 0x06E8
    x"B5",x"76",x"7A",x"32",x"A1",x"77",x"0E",x"00", -- 0x06F0
    x"21",x"80",x"74",x"06",x"01",x"CD",x"68",x"77", -- 0x06F8
    x"DA",x"D6",x"76",x"77",x"2C",x"C2",x"FB",x"76", -- 0x0700
    x"51",x"06",x"01",x"CD",x"68",x"77",x"DA",x"D6", -- 0x0708
    x"76",x"BA",x"C2",x"B5",x"76",x"3A",x"A1",x"77", -- 0x0710
    x"47",x"3A",x"A2",x"77",x"B8",x"CA",x"26",x"77", -- 0x0718
    x"3C",x"B8",x"C2",x"32",x"77",x"C9",x"CD",x"2C", -- 0x0720
    x"77",x"C3",x"9C",x"76",x"3E",x"06",x"CD",x"8B", -- 0x0728
    x"77",x"C9",x"06",x"01",x"CD",x"68",x"77",x"D2", -- 0x0730
    x"32",x"77",x"3E",x"24",x"CD",x"8B",x"77",x"06", -- 0x0738
    x"01",x"CD",x"68",x"77",x"D2",x"3F",x"77",x"3E", -- 0x0740
    x"20",x"CD",x"8B",x"77",x"C3",x"00",x"00",x"3A", -- 0x0748
    x"A2",x"77",x"3C",x"32",x"A2",x"77",x"C9",x"2A", -- 0x0750
    x"A4",x"77",x"EB",x"21",x"80",x"74",x"01",x"80", -- 0x0758
    x"00",x"ED",x"B0",x"EB",x"22",x"A4",x"77",x"C9", -- 0x0760
    x"D5",x"11",x"EE",x"1B",x"DB",x"25",x"E6",x"01", -- 0x0768
    x"C2",x"82",x"77",x"1D",x"C2",x"6C",x"77",x"15", -- 0x0770
    x"C2",x"6C",x"77",x"05",x"C2",x"69",x"77",x"D1", -- 0x0778
    x"37",x"C9",x"DB",x"20",x"D1",x"F5",x"81",x"4F", -- 0x0780
    x"F1",x"B7",x"C9",x"F5",x"DB",x"25",x"E6",x"20", -- 0x0788
    x"CA",x"8C",x"77",x"F1",x"D3",x"20",x"C9",x"AF", -- 0x0790
    x"67",x"6F",x"11",x"00",x"40",x"CD",x"82",x"1F", -- 0x0798
    x"C9",x"00",x"00",x"00",x"00",x"00",x"58",x"4D", -- 0x07A0
    x"4F",x"44",x"45",x"4D",x"28",x"43",x"48",x"45", -- 0x07A8
    x"43",x"4B",x"53",x"55",x"4D",x"29",x"3A",x"33", -- 0x07B0
    x"38",x"34",x"30",x"30",x"2C",x"38",x"2C",x"4E", -- 0x07B8
    x"2C",x"31",x"50",x"52",x"45",x"53",x"53",x"20", -- 0x07C0
    x"27",x"2A",x"27",x"20",x"4F",x"52",x"20",x"27", -- 0x07C8
    x"23",x"27",x"20",x"54",x"4F",x"20",x"44",x"4F", -- 0x07D0
    x"57",x"4E",x"4C",x"4F",x"41",x"44",x"20",x"20", -- 0x07D8
    x"20",x"20",x"44",x"4F",x"57",x"4E",x"4C",x"4F", -- 0x07E0
    x"41",x"44",x"49",x"4E",x"47",x"2E",x"2E",x"2E", -- 0x07E8
    x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20", -- 0x07F0
    x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"FF"  -- 0x07F8
  );


    -- pragma translate_off
    -- := (others => (others => '0'))
    -- pragma translate_on
   

begin

  mem: process (clk_i)
  begin

    if clk_i'event and clk_i = '1' then
      if we_i = '1' then
        mem_q(to_integer(unsigned(a_i))) <= d_i;
      end if;

      d_o <= mem_q(to_integer(unsigned(a_i)));
    end if;

  end process mem;

end rtl;
