// Teclas no extendidas
`define KEY_RELEASED 8'hf0
`define KEY_EXTENDED 8'he0
`define KEY_ESC 	8'h76
`define KEY_F1 		8'h05
`define KEY_F2 		8'h06
`define KEY_F3 		8'h04
`define KEY_F4 		8'h0C
`define KEY_F5 		8'h03
`define KEY_F6 		8'h0B
`define KEY_F7 		8'h83
`define KEY_F8 		8'h0A
`define KEY_F9 		8'h01
`define KEY_F10 	8'h09
`define KEY_F11 	8'h78
`define KEY_F12 	8'h07

`define KEY_BL 		8'h0E
`define KEY_1 		8'h16
`define KEY_2 		8'h1E
`define KEY_3 		8'h26
`define KEY_4 		8'h25
`define KEY_5 		8'h2E
`define KEY_6 		8'h36
`define KEY_7 		8'h3D
`define KEY_8 		8'h3E
`define KEY_9 		8'h46
`define KEY_0 		8'h45
`define KEY_APOS 	8'h4E
`define KEY_AEXC 	8'h55
`define KEY_BKSP 	8'h66

`define KEY_TAB 	8'h0D
`define KEY_Q 		8'h15
`define KEY_W 		8'h1D
`define KEY_E 		8'h24
`define KEY_R 		8'h2D
`define KEY_T 		8'h2C
`define KEY_Y 		8'h35
`define KEY_U 		8'h3C
`define KEY_I 		8'h43
`define KEY_O 		8'h44
`define KEY_P 		8'h4D
`define KEY_CORCHA 	8'h54
`define KEY_CORCHC 	8'h5B
`define KEY_ENTER 	8'h5A

`define KEY_CPSLK 	8'h58
`define KEY_A 		8'h1C
`define KEY_S 		8'h1B
`define KEY_D 		8'h23
`define KEY_F 		8'h2B
`define KEY_G 		8'h34
`define KEY_H 		8'h33
`define KEY_J 		8'h3B
`define KEY_K 		8'h42
`define KEY_L 		8'h4B
`define KEY_NT 		8'h4C
`define KEY_LLAVA 	8'h52
`define KEY_LLAVC 	8'h5D

`define KEY_LSHIFT	8'h12
`define KEY_LT 		8'h61
`define KEY_Z 		8'h1A
`define KEY_X 		8'h22
`define KEY_C 		8'h21
`define KEY_V 		8'h2A
`define KEY_B 		8'h32
`define KEY_N 		8'h31
`define KEY_M 		8'h3A
`define KEY_COMA 	8'h41
`define KEY_PUNTO 	8'h49
`define KEY_MENOS 	8'h4A
`define KEY_RSHIFT	8'h59

`define KEY_LCTRL 	8'h14
`define KEY_LALT 	8'h11
`define KEY_SPACE 	8'h29

`define KEY_KP0 	8'h70
`define KEY_KP1 	8'h69
`define KEY_KP2 	8'h72
`define KEY_KP3 	8'h7A
`define KEY_KP4 	8'h6B
`define KEY_KP5 	8'h73
`define KEY_KP6 	8'h74
`define KEY_KP7 	8'h6C
`define KEY_KP8 	8'h75
`define KEY_KP9 	8'h7D
`define KEY_KPPUNTO 8'h71
`define KEY_KPMAS 	8'h79
`define KEY_KPMENOS 8'h7B
`define KEY_KPASTER 8'h7C

`define KEY_BLKNUM	8'h77
`define KEY_BLKSCR 	8'h7E

// Teclas extendidas (E0 + scancode)
`define KEY_WAKEUP 	8'h5E
`define KEY_SLEEP 	8'h3F
`define KEY_POWER 	8'h37
`define KEY_INS 	8'h70
`define KEY_SUP 	8'h71
`define KEY_HOME 	8'h6C
`define KEY_END 	8'h69
`define KEY_PGU 	8'h7D
`define KEY_PGD 	8'h7A
`define KEY_UP 		8'h75
`define KEY_DOWN 	8'h72
`define KEY_LEFT 	8'h6B
`define KEY_RIGHT 	8'h74
`define KEY_RCTRL 	8'h14
`define KEY_ALTGR 	8'h11
`define KEY_KPENTER 8'h5A
`define KEY_KPSLASH 8'h4A
`define KEY_PRTSCR 	8'h7C
