-------------------------------------------------------------------------------
--
-- Synthesizable model of TI's TMS9918A, TMS9928A, TMS9929A.
--
-- $Id: vdp18_sprite-c.vhd,v 1.3 2006/06/18 10:47:06 arnim Exp $
--
-------------------------------------------------------------------------------

configuration vdp18_sprite_rtl_c0 of vdp18_sprite is

  for rtl
  end for;

end vdp18_sprite_rtl_c0;
