-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity VIC20_CARTRIDGE2 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of VIC20_CARTRIDGE2 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "8808D919DD57155551DB4619661DB4786A79D175D164599618C08118B855B110";
    attribute INIT_01 of inst : label is "2790483658161506D5CA126A7FA405841B524261A000000A2354865230880020";
    attribute INIT_02 of inst : label is "9527572540548E7FAD20D1601D8982F140D93E48E7FAD23F77923C9D8523E43A";
    attribute INIT_03 of inst : label is "01018C7C10E06C48631F041B121177B431E4CC1AC8F9501E4CC38C8C93306B22";
    attribute INIT_04 of inst : label is "411515435750959404802B84845B00005B00005B2000582ECD89058B0817580A";
    attribute INIT_05 of inst : label is "181306432C914320628904174D03241D3408856081179A3495349141D1413491";
    attribute INIT_06 of inst : label is "104437142C22C66ACC5ACD9D471D4D9AB8C4426A3416404CC4C204514056DADA";
    attribute INIT_07 of inst : label is "A004162D5379B15C4950D22841976250B928180AC095174ACCD282E920912C00";
    attribute INIT_08 of inst : label is "8982830046CA4DB080647044D6249044D63A065DC983014B0C17580679B15F48";
    attribute INIT_09 of inst : label is "916CD019501208E9500340654048C9624904245049281145042E141349146DAD";
    attribute INIT_0A of inst : label is "7CAF1927C291CB15C46B54B21355D64287A2B6919615D092E69DA61A579A6986";
    attribute INIT_0B of inst : label is "D715D444CA727008C57111249E4B55D44A9440E88022DA56D5A4744154515B6B";
    attribute INIT_0C of inst : label is "181E02340071019A82091349E054D00952092142440BB164C0815374911D9C40";
    attribute INIT_0D of inst : label is "8861434D8143A0D2E0DF6795D607A468A08DD8D0915D11741A07A22758241998";
    attribute INIT_0E of inst : label is "080951A44545C851209D4D42743417149D23496111174192545425445122340D";
    attribute INIT_0F of inst : label is "2D2086C0A4B0360DD454374141714D50DE3176011C0C950D0958D4104941135B";
    attribute INIT_10 of inst : label is "4DD3741DC20274126805124114D24114D68084926A6474510181E0205903364A";
    attribute INIT_11 of inst : label is "049034121624068205981045355A0181E1995591741535614D42850549991D06";
    attribute INIT_12 of inst : label is "20241014674640607837634D1D022466474534535A0181E10075098075098505";
    attribute INIT_13 of inst : label is "6CC9A04134D0460D3601045D551D0302045340801E407157FA3FA3F0767645D0";
    attribute INIT_14 of inst : label is "6C595B69DB469DB514405876B44744089511816451D0145703B0E415D0919155";
    attribute INIT_15 of inst : label is "16405876B447440815E3281662468955D42078D01556DA46D45D160C116DAD15";
    attribute INIT_16 of inst : label is "A810809014DA8159E42078D01756DA46D455160C916DAD257C515B691B5691B5";
    attribute INIT_17 of inst : label is "2B02C2864C04810320402412493542017B7D81E4E459E2045430830CC0464E06";
    attribute INIT_18 of inst : label is "37624DD10E10C2A7103A46744D9306C2090305089D812750D819CAC598C9424C";
    attribute INIT_19 of inst : label is "4934E30C1B0124C28D534DC144D0D4014D834244C2A2400A1053414D9D28C34A";
    attribute INIT_1A of inst : label is "4D093B04D81B14285060681C0D10D05042090506174248510511AE114445D674";
    attribute INIT_1B of inst : label is "273498860244C0C344C037273490D400230136A845DC9350241302B30489D391";
    attribute INIT_1C of inst : label is "0730065045CD161DAD2E12835483752114138C9CD05CB4C9860244CCC344CC37";
    attribute INIT_1D of inst : label is "E38ED139F2067C8A4404B443640324341C124912A824D9C019455344555555D4";
    attribute INIT_1E of inst : label is "491450410434AB6D02324113620C614070C92449034005064D108318501C3038";
    attribute INIT_1F of inst : label is "423688004D1F3BCA049345241A4C02824180A13005E4500A8A2E800905060024";
    attribute INIT_20 of inst : label is "4232EA6200A25D000220044109511011234AC88C04CAA04004585B469A696631";
    attribute INIT_21 of inst : label is "9283344205504514504C0CA328424D536A18A3976074050656458C0954914CA1";
    attribute INIT_22 of inst : label is "33714D955912965186A83452C611C6112014544482545C0D1061454741681121";
    attribute INIT_23 of inst : label is "20800B01D10E910AA56924D06936939341CA9DA45B3B364F38114452D3235681";
    attribute INIT_24 of inst : label is "244AA001B3447641D091124746C9241D0A38C00924274AA1D098D91373B04801";
    attribute INIT_25 of inst : label is "000000000F0A28BCECECECECECA8A8A8A8A8A8B016AC09212024118E01D50D28";
    attribute INIT_26 of inst : label is "00000061FDF00FC693CAA357B55ED55C2500FFFFFF1515557A9EA4B100E00700";
    attribute INIT_27 of inst : label is "293FFC0FFC33CC0FFC33CC0FFC33CCEFFBEFFBEFFB2FF88BE2EEBB0000000000";
    attribute INIT_28 of inst : label is "007F40D5C007400B4002AD7F5E2E007F5EFF00000075763FFC000068293FFC68";
    attribute INIT_29 of inst : label is "206D3FE209F5FC46F67BFC7159CFFFC9597FE2014EFF88A5DFFF7615CAB45200";
    attribute INIT_2A of inst : label is "7DB1BD9EFF1C5673FFD2565FFD8053BFE22977FF2D8573FE4E14DAD873D9FFFE";
    attribute INIT_2B of inst : label is "159CFFFC9597F8E014EFC88A5DFFF7615CFF938536B61CF67FFFE81B4FF8827D";
    attribute INIT_2C of inst : label is "FC88053BFE22977FDDD8573FFFE14DAD873D9FFFFE06D3FFA09F5FC46F67BFE2";
    attribute INIT_2D of inst : label is "A5DFF93615CFFFF8536B61CF67FFFF8DB4FFF827D7F11BD9EFF885673FFB2565";
    attribute INIT_2E of inst : label is "FFFE14DAD873D9FFFFE26D3FE209F5FC46F67BFF9159CFF6C9597F00014EFC6C";
    attribute INIT_2F of inst : label is "86858C292129212921F246464647C9951D959951D95338D7A3A020B0751E04E7";
    attribute INIT_30 of inst : label is "6C151D1D151511111D1D1D1D15151111111D1D1D15151515151D1515151DBD86";
    attribute INIT_31 of inst : label is "F1F1730547474547454747454747474547474747474747474747474547474745";
    attribute INIT_32 of inst : label is "7C5C7C5C7CC171F1F1717131F1317171F1F17131713171F1F1F17131F1317171";
    attribute INIT_33 of inst : label is "FFFFFFFFFFFFFFF07C5C7C5C7C5C7C5C7C5C7C5C7C5C7C5C7C5C7C5C7C5C7C5C";
    attribute INIT_34 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_35 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_37 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "C00011E561C8761C87A2D8F2E83A3FB80E0C322CB23C8F23CFC8A31AB20F0023";
    attribute INIT_01 of inst : label is "0600083F8C0CBA0C764832D05713C32C31D282C3480000CD3D4A2F880C000000";
    attribute INIT_02 of inst : label is "3297710630108C571020FE323688C4CA06623108C5718231148231D100230670";
    attribute INIT_03 of inst : label is "2320CD5FC1F005081F57F001421097F931720D1748C18C1720D0748D04341923";
    attribute INIT_04 of inst : label is "EF29963D494F5253C32C31EC0020E40820E448E0E408E2C78646C60B4423CC8D";
    attribute INIT_05 of inst : label is "38E0150C28820810300710ADAE2216B6B888AF84AB9CF09E72AEB9E758E3BEFB";
    attribute INIT_06 of inst : label is "38D8091A2D226C8004600A9ECBB0A29A83ECA2663908515B0409A02BC25A5A5E";
    attribute INIT_07 of inst : label is "01F8533B297171C4018C8200C989516255288CC0E2B2ADA0046002C0C73D2D32";
    attribute INIT_08 of inst : label is "88CC43CBC8008A00218F0108930F710893142625851E234B4823CC8CB171C608";
    attribute INIT_09 of inst : label is "324E68018C021BC18C09A0063008C530F7109C91A79E72469E758E3BEFBCA5A5";
    attribute INIT_0A of inst : label is "740D0117409E09B6ECB379520136CCB2A562FBE2EBA21D225D367DB4DB7CFFEF";
    attribute INIT_0B of inst : label is "7DF2FCA4FE92BF0C7CBF2B2A7509B2EEA81486480C99E79BEAFA874BEAF96969";
    attribute INIT_0C of inst : label is "7A7509BAA89709A8004200AB5ACAE22B293290AAC0AD5084E2232BEA32D614A7";
    attribute INIT_0D of inst : label is "84208AEFA30BD2B05CD6F57D4E9D549C4C0DE880DADAD5E57A9D62AF909E3A3A";
    attribute INIT_0E of inst : label is "268D9A40426D84928E3A4D88E8350B1A3D90A319A18F6FDBF6F482409250282B";
    attribute INIT_0F of inst : label is "EEA841849AB89D27AC909EA270B1A79A70C0952B248869A7861CA49AC26F9AC4";
    attribute INIT_10 of inst : label is "A768EAA2C9A8CAA8E42669E39EF8EF8EB8D26868E68A8A66A7A758DC219C1944";
    attribute INIT_11 of inst : label is "AE3A0AB09E9E27CD421C6167BCA3A7A75D252E58F8D68FA3A38DC6348525DA9C";
    attribute INIT_12 of inst : label is "9A8EA099A8A8A9E9D48E92A3DA0D15B976A7BE3AE3A7A7502AE9238AE8234206";
    attribute INIT_13 of inst : label is "404A49EF8EBAC82F9E23AC5651EE2380AE79C892F48AF09421821823596963E4";
    attribute INIT_14 of inst : label is "AF5257DF6FCBFE87BD92FA5696488880250350841EE2169789C274A5F0106149";
    attribute INIT_15 of inst : label is "BC92FA569648888065AC3508634D025D4EA9D6621797FFCA1EFABD206BE5A534";
    attribute INIT_16 of inst : label is "009D10527CDD065D5EA9D6621697FFCA1EFEBD202BE5A534AF5657DF6FDBF687";
    attribute INIT_17 of inst : label is "038CE105ABA70AE8C2F0AE7BE334A28AD35BA758DC210D1A7CBE4BE388C5ABA7";
    attribute INIT_18 of inst : label is "9DB1A71681D0E30529D56945A768E7C4422228027A0A0792BCA5C102188109CE";
    attribute INIT_19 of inst : label is "06BC0C2F9E239CE3232BA389CA7AB809EB88C9C8E3118227D278E9E76F30E3CC";
    attribute INIT_1A of inst : label is "AFC2BF0AFC2B0A3028F2A02F2B28AC68E3868C1A8FC88A3023E83C920E78F0FA";
    attribute INIT_1B of inst : label is "180A384981A6408BE60CBC1B0A3CA989BC23AE5002546BF35453880129232BC1";
    attribute INIT_1C of inst : label is "997CBCA1AF82BE95A590F24BCACBC7401A303064A8F3BA494981A6448BE600BC";
    attribute INIT_1D of inst : label is "BAEB9A163007840FCABEFCAAEA882AAC00414A2AAB16B9F2F2425ACAF25E5D4E";
    attribute INIT_1E of inst : label is "AFBEFBEFBEAE9965AA242F0AE127208AE490AC2390A22BBC2B0049C822B93CAE";
    attribute INIT_1F of inst : label is "A01A4AABEB2D17409EF8EF8EF9884A48AF0A9802A73A7A090995C92927BC2ABC";
    attribute INIT_20 of inst : label is "6A8255598A42258908AA249120909A9293898488BC8AABC2A48810C43A6A5814";
    attribute INIT_21 of inst : label is "69483920C9212940596C099264B10D2B743742723074298A65A9448A809A6991";
    attribute INIT_22 of inst : label is "82908162111244711EA43EB24D32CF3201D49556C82404CE40214954A51011A9";
    attribute INIT_23 of inst : label is "52AA8C231EC11E414DB38E29D38F3BF2A30936CC9025244F38521C1EE92BC902";
    attribute INIT_24 of inst : label is "28AAA5053E77608D80FD23F794F20C583424C8A3082A2AA510E4E232005140C5";
    attribute INIT_25 of inst : label is "40040040040F34DDFECFDCEDFECFDCEDFECFDC0E380086012A2C62402512D983";
    attribute INIT_26 of inst : label is "FF0000069B0690EFFB7FFD6FFC3FF93FE800FFFFFF1E40000E4390AC00500400";
    attribute INIT_27 of inst : label is "FC27D833FC3CFC33FC3CFC33FC3CFC4FF14FF14FF1ABEADFF74FF100000000FF";
    attribute INIT_28 of inst : label is "005540554001E00E000AFDE7AD7900EFADFD000000C245FFFF00003FFC25583F";
    attribute INIT_29 of inst : label is "D41080361002052440B8021080F000020CC00D1C0F00D840CC012483C6475711";
    attribute INIT_2A of inst : label is "827D102E0084203C003083300A0703C0361033003520F300876105392902D000";
    attribute INIT_2B of inst : label is "080F000820CC0F41C0F002C40CC012483CC021D8414E4A40B4000504200D8400";
    attribute INIT_2C of inst : label is "00E0703C0361033013520F300276105392902D000141080021002052440B800D";
    attribute INIT_2D of inst : label is "40CC04D483CC009D8414E4A40B4000584200084008149102E0034203C0060833";
    attribute INIT_2E of inst : label is "00036105392902D000151080361002052440B8009080F001820CC0391C0F0318";
    attribute INIT_2F of inst : label is "80809C050D01090D05F075465767CC840840C840840F85CEF5FD9A041916C557";
    attribute INIT_30 of inst : label is "DC03070B0F03070707070B0B0F0F030303070B0B0F0F0303030B0303030B75C3";
    attribute INIT_31 of inst : label is "A0602B00C1C0C0C1C0C0C1C0C1C0C1C0C1C0C1C1C1C0C1C1C1C0C2C0C1C0C2C0";
    attribute INIT_32 of inst : label is "280828082AC02060A0E02020A02020E0A060202020202060A0602020A02020E0";
    attribute INIT_33 of inst : label is "FFFFFFFFFFFFFFF0280828082808280828082808280828082808280828082808";
    attribute INIT_34 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_35 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_37 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "12B288E8E138466098600800084A01B2606142614260942614ED11127B580C88";
    attribute INIT_01 of inst : label is "90443642BE40064002D018C90048100900B45843200000C9A10901853B2040C8";
    attribute INIT_02 of inst : label is "CE4B009106C36D0040D90AF902D3EEFFE4054136D0040DB6010DB50450DB5044";
    attribute INIT_03 of inst : label is "52DBEC1009091536B30402454D9C9B01480021B036D44180021B036D4586C0D9";
    attribute INIT_04 of inst : label is "1020028101A0002810010003C54903014923614903214082303070BBABA5BE40";
    attribute INIT_05 of inst : label is "A6B87AA8A2BAA8AAFBA8A2409ED8C9027B6D152D155732410241041005144104";
    attribute INIT_06 of inst : label is "241941C1EEB4648B2EE27026699DE2282462848350C287A410D48325C90A202B";
    attribute INIT_07 of inst : label is "EA8DEF9CE4B44802E4410DBAB380BCA44B4D3EE28992649B2E22D9E82C93EE8D";
    attribute INIT_08 of inst : label is "D3EEAA651B22EAC8BBA4CA2D2FA48A2D2F81CE027292521BA3A5BE40B4480036";
    attribute INIT_09 of inst : label is "126C02B4410DACF441A00AD1043672FA48A24486134D12104D3265955554A202";
    attribute INIT_0A of inst : label is "AE2B88CAE20ED192648B014DB592648C8CA4659A5552DC9475D2655449D75955";
    attribute INIT_0B of inst : label is "4102439D488410E54090E4C132D11246909089BB254996499264B77579742880";
    attribute INIT_0C of inst : label is "3132D489657724223212849324496D9106004CA4E344842A8990670902024DD3";
    attribute INIT_0D of inst : label is "76EB64D117D47D32B20CC330CE4C90A2B36823B286828CE3384CB447AA617A79";
    attribute INIT_0E of inst : label is "52946186859634425D56161579D960C9564E1784285D1344D13D05849908C093";
    attribute INIT_0F of inst : label is "22436A5A892264596165679D960C9965B9049BD9236D465B34A30546C91344EB";
    attribute INIT_10 of inst : label is "9826199A94256995D89276176136136139F52745D29D9D2793132D0D0A90C9AA";
    attribute INIT_11 of inst : label is "65A6E1B2606B58F010A9291844A7931320240E663A06618D1AD0D280A4060260";
    attribute INIT_12 of inst : label is "4255B249E9D9E4C4CA618D1A0250903980984D84E793132966585A1679DA5872";
    attribute INIT_13 of inst : label is "B2E6241A41A60A5C6A506A4E64EEDA2261A62D0DB296849800C00C08093998ED";
    attribute INIT_14 of inst : label is "A8406659266996B75425798809088361268C042A4EED901A2605A126B8A52501";
    attribute INIT_15 of inst : label is "542579880908836126A0C0428CA03260CDA4C82D9399966ADD5E5F6125E20280";
    attribute INIT_16 of inst : label is "A17A953DE7203260CDA4C82D9399966ADD5E5F6125E20280A040665926699AB7";
    attribute INIT_17 of inst : label is "9A2288919C1CA707098271C61680B435C8339325050A9261E970371ED4119C9C";
    attribute INIT_18 of inst : label is "4286124654AA899374C9019190A410E632D8C0890212938DE3261450A37694A8";
    attribute INIT_19 of inst : label is "B47A905E48504A899027121409E5E5741E14A40A898D1C92A9049490AB9A8AE6";
    attribute INIT_1A of inst : label is "1E1271C1E361492F448C8F299463030490504ACA4AE6F90850458E426919663B";
    attribute INIT_1B of inst : label is "D2E17B54B5191737197771D0E17904244E504D1A326147AC436A26CBA890279D";
    attribute INIT_1C of inst : label is "4CA6509C97925E620249243709373728C12A410304AC8B3654B5191B37197F71";
    attribute INIT_1D of inst : label is "45140E07DC81FB273951739509D0CB58B28B112800F9429942326519524E60CE";
    attribute INIT_1E of inst : label is "934535914D5B488210985B16CD1BEB66D2616C5244059B64D93B46FAD9B4A651";
    attribute INIT_1F of inst : label is "8C892AA5142B8AE2513513513657D015532A674095CD7D2626325F40554CA944";
    attribute INIT_20 of inst : label is "AAA4AAA8D284AA28220193840161664E0CA6903E4FE004CA92BA0EC3B98108C8";
    attribute INIT_21 of inst : label is "64D8F0C276D8C432082324499B8CB82EA86A86A6DF288A0AA09AD009B28A244A";
    attribute INIT_22 of inst : label is "CD042042202983F0FE1240A44512451A2080880990587E3C32E8088092210246";
    attribute INIT_23 of inst : label is "82AA40D28E188E58749D49241F41F79412D1D2749B43CB2DBA826AC22CC449A2";
    attribute INIT_24 of inst : label is "44A00D2FC35B7BE4E904E490BF0FB2DEBC7E12ACBE47A00FD3CBCF9FA76FCADA";
    attribute INIT_25 of inst : label is "00000000000518564764764754754754654654C3B8B2E22B4044D2229DD2DDFC";
    attribute INIT_26 of inst : label is "FF096700000960BFFEDFF79FFC3FF61D6000FFFFFF8040001004000000200000";
    attribute INIT_27 of inst : label is "FF41413CFC3F3C3CFC3F3C3CFC3F3CEFFBEFFBEFFB7FFD8FF2EFFB0000FFFFFF";
    attribute INIT_28 of inst : label is "80D5406DC00D4001E00BF4FFFA7F00FFFE7C0096001400FFFF0000FFFF0000FF";
    attribute INIT_29 of inst : label is "C3042AAF0C10AA952072AA9481CAAA83002AA5401CAABC2002AA94C0DEDFEC95";
    attribute INIT_2A of inst : label is "2A95481CAAA52072AAB0C00AA550072AAF0800AA953037AABF3042954081CAAB";
    attribute INIT_2B of inst : label is "481CAAAC3002A55401CABFC2002AA94C0DEAAFCC10A5502072AAB0C10AABC304";
    attribute INIT_2C of inst : label is "AA550072AAF0800AA953037AAAF3042954081CAAA82042AAF0C10AA952072AA5";
    attribute INIT_2D of inst : label is "2002AA54C0DEAABCC10A5502072AAA0410AAAC3042AA5481CAA952072AAF0C00";
    attribute INIT_2E of inst : label is "AAAB3042954081CAAA81042AAF0C10AA952072AA5481CAAFC3002A95401CAAFC";
    attribute INIT_2F of inst : label is "01021C080404000C0CB001223303CCCCC888CCCC888BA75229392E0000000003";
    attribute INIT_30 of inst : label is "1C0404040408080804040404040400000004040404040404040404040404BFC3";
    attribute INIT_31 of inst : label is "40404B0101000101010001010100010101000101010001010300010103000101";
    attribute INIT_32 of inst : label is "1020102011C04040404080004000804040404000400040404040400040008040";
    attribute INIT_33 of inst : label is "FFFFFFFFFFFFFFF0102010201020102010201020102010201020102010201020";
    attribute INIT_34 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_35 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_37 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "22A8222220A82A89A22288A288AE2BB88B8A2A8A268BA2A8A26FC22BB98BF188";
    attribute INIT_01 of inst : label is "15542C89A088228822CC2B895559620A20B33BC2200000C2A4892884228008A0";
    attribute INIT_02 of inst : label is "610B55155402CD5550B2268022FECAC00555542CD5550B34550B355550B35555";
    attribute INIT_03 of inst : label is "C292CD555151542CB75554550B0C0B55515545042CD55515545042CD551410B0";
    attribute INIT_04 of inst : label is "8222229484A52129620A20B333396333B97333397333B0827B7B7BFBC708A00C";
    attribute INIT_05 of inst : label is "28B0CA082C82882CB28A2C0A4090C829024CC22CC20A22082208208220820820";
    attribute INIT_06 of inst : label is "2088CCECEF33B88A8AE2232388E8A0296938808CCCCC9CA533F3F300888A1028";
    attribute INIT_07 of inst : label is "A21F2B0E10B5515405550B2832848C9CCBFFAC228022098A8AE2A2E865B7EF0C";
    attribute INIT_08 of inst : label is "FEC2B2408A82A6A0ABADA2CF2B2DA2CF2B08CA123287C23BC308AC08B551542C";
    attribute INIT_09 of inst : label is "662D5405552B2DC55505501554AC3282DA2C0889C20C2223083208208208A102";
    attribute INIT_0A of inst : label is "AC2B08CAC222CEE2398B552B3EA2298F88B31862186688B39AE29A6988638618";
    attribute INIT_0B of inst : label is "BAE2384F3CC8CE23B88E108C22CEE2394888802E8F3E69886619A230B0222840";
    attribute INIT_0C of inst : label is "1022F384B1AA222232304C02209409020A518C20930C8CC98086208822222A82";
    attribute INIT_0D of inst : label is "3B92418646F1F062B52A8AA2AA0888A4A6C2202222262A8AA808BF1BA9386AA8";
    attribute INIT_0E of inst : label is "CFF32CC88842232218620231B8088C04611DC62222188621886C888988888C86";
    attribute INIT_0F of inst : label is "6123B2B384A008C220230B8088C042102A4C08C2233231027B2637308886218A";
    attribute INIT_10 of inst : label is "8E2398E6F3F198E1888AA386386386386ABCF6318AA4A8AA8102273732A4C09B";
    attribute INIT_11 of inst : label is "38D0DCE23938CF333327048E18AA810222220C23B926398DCE33304892022638";
    attribute INIT_12 of inst : label is "3F18E22AAA4AA04089398DCE26334830898E18E1AA810227F3880E33B80E2301";
    attribute INIT_13 of inst : label is "A8AE2182182088C308C7092C2210920208A09CCCA2308C081041041488B08EEF";
    attribute INIT_14 of inst : label is "A92029A6219866A2080C284408841E47024CCCC92109084A00CC3302808CCC80";
    attribute INIT_15 of inst : label is "080C284408841E470294CCCC8C913022A46089090B08618A882C0BF300A10248";
    attribute INIT_16 of inst : label is "630D8CCC27213022A46089090B08618A882C0BF300A10248A52029A6219866A2";
    attribute INIT_17 of inst : label is "0A02808A82C260B0882208208E48B33388AA82233332A4DC230F30C231CA82C2";
    attribute INIT_18 of inst : label is "198DC62233B1808AA0888488866086E23090CC8862324B8CA302333320327198";
    attribute INIT_19 of inst : label is "2309A4C318C7198082134231CC90A331CA0091898088CCC6B060418668098202";
    attribute INIT_1A of inst : label is "C2320CCC2308C872318C232902233331876318C20A02F824C3962E0888822899";
    attribute INIT_1B of inst : label is "8CDC63F3F8C42630C4270C8DDC62322219C718A9302230A9332602A2A88220CC";
    attribute INIT_1C of inst : label is "08A4088C02F00A11022A7330C430E224CC66923231A98C32F3F8C42230C4230C";
    attribute INIT_1D of inst : label is "0000260B8A00E283840A384084FC0C08A8B0A22954C8229022302098222C22AA";
    attribute INIT_1E of inst : label is "42081082040B28426648822088C29240892208810DCCC208822230A490226400";
    attribute INIT_1F of inst : label is "8CC89990822B0AC2082082082220CB30C22F2FCFC2842C222232232CC308BF08";
    attribute INIT_20 of inst : label is "A67F0001F8C8C2222266488CF22211224C12F3E00A05508BC8A42B8AE84888CC";
    attribute INIT_21 of inst : label is "22FCFCB20290B222249F22248A93E2308CCCCCC88C0892448842F3C222249224";
    attribute INIT_22 of inst : label is "09C9D28022248AA2AA0988BF8A22082220484886FC88A43F2290848842322113";
    attribute INIT_23 of inst : label is "35990CC222332233B88E0461AE18E08CC6CEE23988CCCA0E3C2289A630E18A97";
    attribute INIT_24 of inst : label is "88A5522284888A022620C8880A1824224CCDF3F92088A55227F3F81C8CCC89F2";
    attribute INIT_25 of inst : label is "00000000010000033222111000333222111000A698A8A2273A88222252222261";
    attribute INIT_26 of inst : label is "FF92FE0000F00FC553C963AB7AADEA540500FFFFFF0000000000015400100100";
    attribute INIT_27 of inst : label is "FF00000FFC33FC0FFC33FC0FFC33FC4FF14FF14551FFFFDD7747D1FFFFFFFFFF";
    attribute INIT_28 of inst : label is "405540554007800B407FF0FFFF7FE0FFFF1E406067000015540000FFFF0000FF";
    attribute INIT_29 of inst : label is "C004157F041050000071540001C55540041540041C55FC1041540041CB9A8A55";
    attribute INIT_2A of inst : label is "1400001C5500007155700105500107157F04105500107357FF0040000001C557";
    attribute INIT_2B of inst : label is "001C555C0041500041C57FC1041540041CD5FFC01000000071557001055FC104";
    attribute INIT_2C of inst : label is "5400107157F041054001073557F0040000001C5554004155F041050000071540";
    attribute INIT_2D of inst : label is "1041500041CD55FC010000000715550010555C1041400001C5500007155F0010";
    attribute INIT_2E of inst : label is "55570040000001C5554004157F041050000071550001C55FC0041500041C57FC";
    attribute INIT_2F of inst : label is "03030C8C8C8C8C88883222222230CCCCCCCCCCCCCCC300004120000000000003";
    attribute INIT_30 of inst : label is "0C0C0C0C0C0C0C0C0C0C0C0C0C0C0000000C0C0C0C0C0C0C0C0C0C0C0C0C3BC2";
    attribute INIT_31 of inst : label is "C0C0C30303030303030303030303030303030303030303030203030302030303";
    attribute INIT_32 of inst : label is "3030303030C0C0C0C0C0C000C000C0C0C0C0C000C000C0C0C0C0C000C000C0C0";
    attribute INIT_33 of inst : label is "FFFFFFFFFFFFFFF0303030303030303030303030303030303030303030303030";
    attribute INIT_34 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_35 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_37 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
