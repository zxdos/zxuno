library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package TIA_NTSCLookups is

   constant sync_level: unsigned(7 downto 0) := X"05";
   constant blank_level: unsigned(7 downto 0) := X"5a";

   type lum_lut_type is array (0 to 7) of unsigned(7 downto 0);
   constant lum_lut: lum_lut_type := (
      X"6a",
      X"74",
      X"7e",
      X"88",
      X"91",
      X"9b",
      X"a5",
      X"af");

   type col_lut_type is array (0 to 255) of unsigned(7 downto 0);
   constant col_lut: col_lut_type := (
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"00",
      X"f8",
      X"f1",
      X"ec",
      X"eb",
      X"ec",
      X"f1",
      X"f8",
      X"00",
      X"08",
      X"0f",
      X"14",
      X"15",
      X"14",
      X"0f",
      X"08",
      X"0a",
      X"02",
      X"f9",
      X"f2",
      X"ed",
      X"eb",
      X"ec",
      X"f0",
      X"f6",
      X"fe",
      X"07",
      X"0e",
      X"13",
      X"15",
      X"14",
      X"10",
      X"11",
      X"0b",
      X"03",
      X"fb",
      X"f4",
      X"ee",
      X"eb",
      X"eb",
      X"ef",
      X"f5",
      X"fd",
      X"05",
      X"0c",
      X"12",
      X"15",
      X"15",
      X"15",
      X"12",
      X"0d",
      X"05",
      X"fd",
      X"f5",
      X"ef",
      X"eb",
      X"eb",
      X"ee",
      X"f3",
      X"fb",
      X"03",
      X"0b",
      X"11",
      X"15",
      X"14",
      X"15",
      X"13",
      X"0e",
      X"07",
      X"fe",
      X"f6",
      X"f0",
      X"ec",
      X"eb",
      X"ed",
      X"f2",
      X"f9",
      X"02",
      X"0a",
      X"10",
      X"0f",
      X"14",
      X"15",
      X"14",
      X"0f",
      X"08",
      X"00",
      X"f8",
      X"f1",
      X"ec",
      X"eb",
      X"ec",
      X"f1",
      X"f8",
      X"00",
      X"08",
      X"06",
      X"0e",
      X"13",
      X"15",
      X"14",
      X"10",
      X"0a",
      X"02",
      X"fa",
      X"f2",
      X"ed",
      X"eb",
      X"ec",
      X"f0",
      X"f6",
      X"fe",
      X"fd",
      X"05",
      X"0c",
      X"12",
      X"15",
      X"15",
      X"11",
      X"0b",
      X"03",
      X"fb",
      X"f4",
      X"ee",
      X"eb",
      X"eb",
      X"ef",
      X"f5",
      X"f3",
      X"fb",
      X"03",
      X"0b",
      X"11",
      X"15",
      X"15",
      X"12",
      X"0d",
      X"05",
      X"fd",
      X"f5",
      X"ef",
      X"eb",
      X"eb",
      X"ee",
      X"ed",
      X"f2",
      X"f9",
      X"01",
      X"09",
      X"10",
      X"14",
      X"15",
      X"13",
      X"0e",
      X"07",
      X"ff",
      X"f7",
      X"f0",
      X"ec",
      X"eb",
      X"eb",
      X"ec",
      X"f1",
      X"f8",
      X"00",
      X"08",
      X"0f",
      X"14",
      X"15",
      X"14",
      X"0f",
      X"08",
      X"00",
      X"f8",
      X"f1",
      X"ec",
      X"ed",
      X"eb",
      X"ec",
      X"f0",
      X"f6",
      X"fe",
      X"06",
      X"0e",
      X"13",
      X"15",
      X"14",
      X"10",
      X"0a",
      X"02",
      X"fa",
      X"f2",
      X"f4",
      X"ee",
      X"eb",
      X"eb",
      X"ef",
      X"f5",
      X"fc",
      X"05",
      X"0c",
      X"12",
      X"15",
      X"15",
      X"11",
      X"0b",
      X"04",
      X"fb",
      X"fd",
      X"f5",
      X"ef",
      X"eb",
      X"eb",
      X"ee",
      X"f3",
      X"fb",
      X"03",
      X"0b",
      X"11",
      X"15",
      X"15",
      X"12",
      X"0d",
      X"05",
      X"07",
      X"ff",
      X"f7",
      X"f0",
      X"ec",
      X"eb",
      X"ed",
      X"f2",
      X"f9",
      X"01",
      X"09",
      X"10",
      X"14",
      X"15",
      X"13",
      X"0e");

end TIA_NTSCLookups;

package body TIA_NTSCLookups is

end TIA_NTSCLookups;
