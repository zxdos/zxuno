-------------------------------------------------------------------------------
--
-- FPGA Colecovision
--
-- $Id: cv_bus_mux-c.vhd,v 1.2 2006/01/05 22:25:25 arnim Exp $
--
-------------------------------------------------------------------------------

configuration cv_bus_mux_rtl_c0 of cv_bus_mux is

  for rtl
  end for;

end cv_bus_mux_rtl_c0;
