-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80e3",
     9 => x"f0080b0b",
    10 => x"80e3f408",
    11 => x"0b0b80e3",
    12 => x"f8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"e3f80c0b",
    16 => x"0b80e3f4",
    17 => x"0c0b0b80",
    18 => x"e3f00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80de98",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80e3f070",
    57 => x"80eea827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51b192",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80e4",
    65 => x"800c9f0b",
    66 => x"80e4840c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"e48408ff",
    70 => x"0580e484",
    71 => x"0c80e484",
    72 => x"088025e8",
    73 => x"3880e480",
    74 => x"08ff0580",
    75 => x"e4800c80",
    76 => x"e4800880",
    77 => x"25d03880",
    78 => x"0b80e484",
    79 => x"0c800b80",
    80 => x"e4800c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80e48008",
   100 => x"25913882",
   101 => x"c82d80e4",
   102 => x"8008ff05",
   103 => x"80e4800c",
   104 => x"838a0480",
   105 => x"e4800880",
   106 => x"e4840853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80e48008",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"e4840881",
   116 => x"0580e484",
   117 => x"0c80e484",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80e484",
   121 => x"0c80e480",
   122 => x"08810580",
   123 => x"e4800c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480e4",
   128 => x"84088105",
   129 => x"80e4840c",
   130 => x"80e48408",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80e484",
   134 => x"0c80e480",
   135 => x"08810580",
   136 => x"e4800c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"e4880cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"e4880c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280e4",
   177 => x"88088407",
   178 => x"80e4880c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80e0",
   183 => x"dc0c8171",
   184 => x"2bff05f6",
   185 => x"880cfdfc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80e488",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80e3",
   208 => x"f00c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"a00bec0c",
  1093 => x"86c72d86",
  1094 => x"c72d86c7",
  1095 => x"2d86c72d",
  1096 => x"86c72d86",
  1097 => x"c72d86c7",
  1098 => x"2d86c72d",
  1099 => x"86c72d86",
  1100 => x"c72d86c7",
  1101 => x"2d86c72d",
  1102 => x"86c72d86",
  1103 => x"c72d86c7",
  1104 => x"2d86c72d",
  1105 => x"86c72d86",
  1106 => x"c72d86c7",
  1107 => x"2d86c72d",
  1108 => x"86c72d86",
  1109 => x"c72d86c7",
  1110 => x"2d86c72d",
  1111 => x"86c72d86",
  1112 => x"c72d86c7",
  1113 => x"2d86c72d",
  1114 => x"86c72d86",
  1115 => x"c72d86c7",
  1116 => x"2d86c72d",
  1117 => x"86c72d86",
  1118 => x"c72d86c7",
  1119 => x"2d86c72d",
  1120 => x"86c72d86",
  1121 => x"c72d86c7",
  1122 => x"2d86c72d",
  1123 => x"86c72d86",
  1124 => x"c72d86c7",
  1125 => x"2d86c72d",
  1126 => x"86c72d86",
  1127 => x"c72d86c7",
  1128 => x"2d86c72d",
  1129 => x"86c72d86",
  1130 => x"c72d86c7",
  1131 => x"2d86c72d",
  1132 => x"86c72d86",
  1133 => x"c72d86c7",
  1134 => x"2d86c72d",
  1135 => x"86c72d86",
  1136 => x"c72d86c7",
  1137 => x"2d86c72d",
  1138 => x"86c72d86",
  1139 => x"c72d86c7",
  1140 => x"2d86c72d",
  1141 => x"86c72d86",
  1142 => x"c72d86c7",
  1143 => x"2d86c72d",
  1144 => x"86c72d86",
  1145 => x"c72d86c7",
  1146 => x"2d86c72d",
  1147 => x"86c72d86",
  1148 => x"c72d86c7",
  1149 => x"2d86c72d",
  1150 => x"86c72d86",
  1151 => x"c72d86c7",
  1152 => x"2d86c72d",
  1153 => x"86c72d86",
  1154 => x"c72d86c7",
  1155 => x"2d86c72d",
  1156 => x"86c72d86",
  1157 => x"c72d86c7",
  1158 => x"2d86c72d",
  1159 => x"86c72d86",
  1160 => x"c72d86c7",
  1161 => x"2d86c72d",
  1162 => x"86c72d86",
  1163 => x"c72d86c7",
  1164 => x"2d86c72d",
  1165 => x"86c72d86",
  1166 => x"c72d86c7",
  1167 => x"2d86c72d",
  1168 => x"86c72d86",
  1169 => x"c72d86c7",
  1170 => x"2d86c72d",
  1171 => x"86c72d86",
  1172 => x"c72d86c7",
  1173 => x"2d86c72d",
  1174 => x"86c72d86",
  1175 => x"c72d86c7",
  1176 => x"2d86c72d",
  1177 => x"86c72d86",
  1178 => x"c72d86c7",
  1179 => x"2d86c72d",
  1180 => x"86c72d86",
  1181 => x"c72d86c7",
  1182 => x"2d86c72d",
  1183 => x"86c72d86",
  1184 => x"c72d86c7",
  1185 => x"2d86c72d",
  1186 => x"86c72d86",
  1187 => x"c72d86c7",
  1188 => x"2d86c72d",
  1189 => x"86c72d86",
  1190 => x"c72d86c7",
  1191 => x"2d86c72d",
  1192 => x"86c72d86",
  1193 => x"c72d86c7",
  1194 => x"2d86c72d",
  1195 => x"86c72d86",
  1196 => x"c72d86c7",
  1197 => x"2d86c72d",
  1198 => x"86c72d86",
  1199 => x"c72d86c7",
  1200 => x"2d86c72d",
  1201 => x"86c72d86",
  1202 => x"c72d86c7",
  1203 => x"2d86c72d",
  1204 => x"86c72d86",
  1205 => x"c72d86c7",
  1206 => x"2d86c72d",
  1207 => x"86c72d86",
  1208 => x"c72d86c7",
  1209 => x"2d86c72d",
  1210 => x"86c72d86",
  1211 => x"c72d86c7",
  1212 => x"2d86c72d",
  1213 => x"86c72d86",
  1214 => x"c72d86c7",
  1215 => x"2d86c72d",
  1216 => x"86c72d86",
  1217 => x"c72d86c7",
  1218 => x"2d86c72d",
  1219 => x"86c72d86",
  1220 => x"c72d86c7",
  1221 => x"2d86c72d",
  1222 => x"86c72d86",
  1223 => x"c72d86c7",
  1224 => x"2d86c72d",
  1225 => x"86c72d86",
  1226 => x"c72d86c7",
  1227 => x"2d86c72d",
  1228 => x"86c72d86",
  1229 => x"c72d86c7",
  1230 => x"2d86c72d",
  1231 => x"86c72d86",
  1232 => x"c72d86c7",
  1233 => x"2d86c72d",
  1234 => x"86c72d86",
  1235 => x"c72d86c7",
  1236 => x"2d86c72d",
  1237 => x"86c72d86",
  1238 => x"c72d86c7",
  1239 => x"2d86c72d",
  1240 => x"86c72d86",
  1241 => x"c72d86c7",
  1242 => x"2d86c72d",
  1243 => x"86c72d86",
  1244 => x"c72d86c7",
  1245 => x"2d86c72d",
  1246 => x"86c72d86",
  1247 => x"c72d86c7",
  1248 => x"2d86c72d",
  1249 => x"86c72d86",
  1250 => x"c72d86c7",
  1251 => x"2d86c72d",
  1252 => x"86c72d86",
  1253 => x"c72d86c7",
  1254 => x"2d86c72d",
  1255 => x"86c72d86",
  1256 => x"c72d86c7",
  1257 => x"2d86c72d",
  1258 => x"86c72d86",
  1259 => x"c72d86c7",
  1260 => x"2d86c72d",
  1261 => x"86c72d86",
  1262 => x"c72d86c7",
  1263 => x"2d86c72d",
  1264 => x"86c72d86",
  1265 => x"c72d86c7",
  1266 => x"2d86c72d",
  1267 => x"86c72d86",
  1268 => x"c72d86c7",
  1269 => x"2d86c72d",
  1270 => x"86c72d86",
  1271 => x"c72d86c7",
  1272 => x"2d86c72d",
  1273 => x"86c72d86",
  1274 => x"c72d86c7",
  1275 => x"2d86c72d",
  1276 => x"86c72d86",
  1277 => x"c72d86c7",
  1278 => x"2d86c72d",
  1279 => x"86c72d86",
  1280 => x"c72d86c7",
  1281 => x"2d86c72d",
  1282 => x"86c72d86",
  1283 => x"c72d86c7",
  1284 => x"2d86c72d",
  1285 => x"86c72d86",
  1286 => x"c72d86c7",
  1287 => x"2d86c72d",
  1288 => x"86c72d86",
  1289 => x"c72d86c7",
  1290 => x"2d86c72d",
  1291 => x"86c72d86",
  1292 => x"c72d86c7",
  1293 => x"2d86c72d",
  1294 => x"86c72d86",
  1295 => x"c72d86c7",
  1296 => x"2d86c72d",
  1297 => x"86c72d86",
  1298 => x"c72d86c7",
  1299 => x"2d86c72d",
  1300 => x"86c72d86",
  1301 => x"c72d86c7",
  1302 => x"2d86c72d",
  1303 => x"86c72d86",
  1304 => x"c72d86c7",
  1305 => x"2d86c72d",
  1306 => x"86c72d86",
  1307 => x"c72d86c7",
  1308 => x"2d86c72d",
  1309 => x"86c72d86",
  1310 => x"c72d86c7",
  1311 => x"2d86c72d",
  1312 => x"86c72d86",
  1313 => x"c72d86c7",
  1314 => x"2d86c72d",
  1315 => x"86c72d86",
  1316 => x"c72d86c7",
  1317 => x"2d86c72d",
  1318 => x"86c72d86",
  1319 => x"c72d86c7",
  1320 => x"2d86c72d",
  1321 => x"86c72d86",
  1322 => x"c72d86c7",
  1323 => x"2d86c72d",
  1324 => x"86c72d86",
  1325 => x"c72d86c7",
  1326 => x"2d86c72d",
  1327 => x"86c72d86",
  1328 => x"c72d86c7",
  1329 => x"2d86c72d",
  1330 => x"86c72d86",
  1331 => x"c72d86c7",
  1332 => x"2d86c72d",
  1333 => x"86c72d86",
  1334 => x"c72d86c7",
  1335 => x"2d86c72d",
  1336 => x"86c72d86",
  1337 => x"c72d86c7",
  1338 => x"2d86c72d",
  1339 => x"86c72d86",
  1340 => x"c72d86c7",
  1341 => x"2d86c72d",
  1342 => x"86c72d86",
  1343 => x"c72d86c7",
  1344 => x"2d86c72d",
  1345 => x"86c72d86",
  1346 => x"c72d86c7",
  1347 => x"2d86c72d",
  1348 => x"86c72d86",
  1349 => x"c72d86c7",
  1350 => x"2d86c72d",
  1351 => x"86c72d86",
  1352 => x"c72d86c7",
  1353 => x"2d86c72d",
  1354 => x"86c72d86",
  1355 => x"c72d86c7",
  1356 => x"2d86c72d",
  1357 => x"86c72d86",
  1358 => x"c72d86c7",
  1359 => x"2d86c72d",
  1360 => x"86c72d86",
  1361 => x"c72d86c7",
  1362 => x"2d86c72d",
  1363 => x"86c72d86",
  1364 => x"c72d86c7",
  1365 => x"2d86c72d",
  1366 => x"86c72d86",
  1367 => x"c72d86c7",
  1368 => x"2d86c72d",
  1369 => x"86c72d86",
  1370 => x"c72d86c7",
  1371 => x"2d86c72d",
  1372 => x"86c72d86",
  1373 => x"c72d86c7",
  1374 => x"2d86c72d",
  1375 => x"86c72d86",
  1376 => x"c72d86c7",
  1377 => x"2d86c72d",
  1378 => x"86c72d86",
  1379 => x"c72d86c7",
  1380 => x"2d86c72d",
  1381 => x"86c72d86",
  1382 => x"c72d86c7",
  1383 => x"2d86c72d",
  1384 => x"86c72d86",
  1385 => x"c72d86c7",
  1386 => x"2d86c72d",
  1387 => x"86c72d86",
  1388 => x"c72d86c7",
  1389 => x"2d86c72d",
  1390 => x"86c72d86",
  1391 => x"c72d86c7",
  1392 => x"2d86c72d",
  1393 => x"86c72d86",
  1394 => x"c72d86c7",
  1395 => x"2d86c72d",
  1396 => x"86c72d86",
  1397 => x"c72d86c7",
  1398 => x"2d86c72d",
  1399 => x"86c72d86",
  1400 => x"c72d86c7",
  1401 => x"2d86c72d",
  1402 => x"86c72d86",
  1403 => x"c72d86c7",
  1404 => x"2d86c72d",
  1405 => x"86c72d86",
  1406 => x"c72d86c7",
  1407 => x"2d86c72d",
  1408 => x"86c72d86",
  1409 => x"c72d86c7",
  1410 => x"2d86c72d",
  1411 => x"86c72d86",
  1412 => x"c72d86c7",
  1413 => x"2d86c72d",
  1414 => x"86c72d86",
  1415 => x"c72d86c7",
  1416 => x"2d86c72d",
  1417 => x"86c72d86",
  1418 => x"c72d86c7",
  1419 => x"2d86c72d",
  1420 => x"86c72d86",
  1421 => x"c72d86c7",
  1422 => x"2d86c72d",
  1423 => x"86c72d86",
  1424 => x"c72d86c7",
  1425 => x"2d86c72d",
  1426 => x"86c72d86",
  1427 => x"c72d86c7",
  1428 => x"2d86c72d",
  1429 => x"86c72d86",
  1430 => x"c72d86c7",
  1431 => x"2d86c72d",
  1432 => x"86c72d86",
  1433 => x"c72d86c7",
  1434 => x"2d86c72d",
  1435 => x"86c72d86",
  1436 => x"c72d86c7",
  1437 => x"2d86c72d",
  1438 => x"86c72d86",
  1439 => x"c72d86c7",
  1440 => x"2d86c72d",
  1441 => x"86c72d86",
  1442 => x"c72d86c7",
  1443 => x"2d86c72d",
  1444 => x"86c72d86",
  1445 => x"c72d86c7",
  1446 => x"2d86c72d",
  1447 => x"86c72d86",
  1448 => x"c72d86c7",
  1449 => x"2d86c72d",
  1450 => x"86c72d86",
  1451 => x"c72d86c7",
  1452 => x"2d86c72d",
  1453 => x"86c72d86",
  1454 => x"c72d86c7",
  1455 => x"2d86c72d",
  1456 => x"86c72d86",
  1457 => x"c72d86c7",
  1458 => x"2d86c72d",
  1459 => x"86c72d86",
  1460 => x"c72d86c7",
  1461 => x"2d86c72d",
  1462 => x"86c72d86",
  1463 => x"c72d86c7",
  1464 => x"2d86c72d",
  1465 => x"86c72d86",
  1466 => x"c72d86c7",
  1467 => x"2d86c72d",
  1468 => x"86c72d86",
  1469 => x"c72d86c7",
  1470 => x"2d86c72d",
  1471 => x"86c72d86",
  1472 => x"c72d86c7",
  1473 => x"2d86c72d",
  1474 => x"86c72d86",
  1475 => x"c72d86c7",
  1476 => x"2d86c72d",
  1477 => x"86c72d86",
  1478 => x"c72d86c7",
  1479 => x"2d86c72d",
  1480 => x"86c72d86",
  1481 => x"c72d86c7",
  1482 => x"2d86c72d",
  1483 => x"86c72d86",
  1484 => x"c72d86c7",
  1485 => x"2d86c72d",
  1486 => x"86c72d86",
  1487 => x"c72d86c7",
  1488 => x"2d86c72d",
  1489 => x"86c72d86",
  1490 => x"c72d86c7",
  1491 => x"2d86c72d",
  1492 => x"86c72d86",
  1493 => x"c72d86c7",
  1494 => x"2d86c72d",
  1495 => x"86c72d86",
  1496 => x"c72d86c7",
  1497 => x"2d86c72d",
  1498 => x"86c72d86",
  1499 => x"c72d86c7",
  1500 => x"2d86c72d",
  1501 => x"86c72d86",
  1502 => x"c72d86c7",
  1503 => x"2d86c72d",
  1504 => x"86c72d86",
  1505 => x"c72d86c7",
  1506 => x"2d86c72d",
  1507 => x"86c72d86",
  1508 => x"c72d86c7",
  1509 => x"2d86c72d",
  1510 => x"86c72d86",
  1511 => x"c72d86c7",
  1512 => x"2d86c72d",
  1513 => x"86c72d86",
  1514 => x"c72d86c7",
  1515 => x"2d86c72d",
  1516 => x"86c72d86",
  1517 => x"c72d86c7",
  1518 => x"2d86c72d",
  1519 => x"86c72d86",
  1520 => x"c72d86c7",
  1521 => x"2d86c72d",
  1522 => x"86c72d86",
  1523 => x"c72d86c7",
  1524 => x"2d86c72d",
  1525 => x"0402dc05",
  1526 => x"0d8059a2",
  1527 => x"902d810b",
  1528 => x"ec0c7a52",
  1529 => x"80e48c51",
  1530 => x"80d4e32d",
  1531 => x"80e3f008",
  1532 => x"792e80f7",
  1533 => x"3880e490",
  1534 => x"0870f80c",
  1535 => x"79ff1256",
  1536 => x"59557379",
  1537 => x"2e8b3881",
  1538 => x"1874812a",
  1539 => x"555873f7",
  1540 => x"38f71858",
  1541 => x"81598075",
  1542 => x"2580d038",
  1543 => x"77527351",
  1544 => x"84a82d80",
  1545 => x"e4e05280",
  1546 => x"e48c5180",
  1547 => x"d7b92d80",
  1548 => x"e3f00880",
  1549 => x"2e9b3880",
  1550 => x"e4e05783",
  1551 => x"fc567670",
  1552 => x"84055808",
  1553 => x"e80cfc16",
  1554 => x"56758025",
  1555 => x"f138b0d9",
  1556 => x"0480e3f0",
  1557 => x"08598480",
  1558 => x"5580e48c",
  1559 => x"5180d788",
  1560 => x"2dfc8015",
  1561 => x"81155555",
  1562 => x"b0960484",
  1563 => x"0bec0c78",
  1564 => x"802e8e38",
  1565 => x"80e0e051",
  1566 => x"b8c72db6",
  1567 => x"ba2db188",
  1568 => x"0480e1c0",
  1569 => x"51b8c72d",
  1570 => x"7880e3f0",
  1571 => x"0c02a405",
  1572 => x"0d0402f0",
  1573 => x"050d840b",
  1574 => x"ec0cb684",
  1575 => x"2db2b92d",
  1576 => x"81f92d83",
  1577 => x"52b5e72d",
  1578 => x"8151858d",
  1579 => x"2dff1252",
  1580 => x"718025f1",
  1581 => x"38840bec",
  1582 => x"0c80df90",
  1583 => x"5186a02d",
  1584 => x"80cb832d",
  1585 => x"80e3f008",
  1586 => x"802e80d6",
  1587 => x"38afd551",
  1588 => x"80de902d",
  1589 => x"80e0e051",
  1590 => x"b8c72db6",
  1591 => x"a62db2c5",
  1592 => x"2db8da2d",
  1593 => x"80e0f40b",
  1594 => x"80f52d80",
  1595 => x"e2ac0870",
  1596 => x"81065455",
  1597 => x"5371802e",
  1598 => x"85387281",
  1599 => x"07537381",
  1600 => x"2a708106",
  1601 => x"51527180",
  1602 => x"2e853872",
  1603 => x"82075372",
  1604 => x"fc0c8652",
  1605 => x"80e3f008",
  1606 => x"83388452",
  1607 => x"71ec0cb1",
  1608 => x"de04800b",
  1609 => x"80e3f00c",
  1610 => x"0290050d",
  1611 => x"0471980c",
  1612 => x"04ffb008",
  1613 => x"80e3f00c",
  1614 => x"04810bff",
  1615 => x"b00c0480",
  1616 => x"0bffb00c",
  1617 => x"0402f405",
  1618 => x"0db3d304",
  1619 => x"80e3f008",
  1620 => x"81f02e09",
  1621 => x"81068a38",
  1622 => x"810b80e2",
  1623 => x"a40cb3d3",
  1624 => x"0480e3f0",
  1625 => x"0881e02e",
  1626 => x"0981068a",
  1627 => x"38810b80",
  1628 => x"e2a80cb3",
  1629 => x"d30480e3",
  1630 => x"f0085280",
  1631 => x"e2a80880",
  1632 => x"2e893880",
  1633 => x"e3f00881",
  1634 => x"80055271",
  1635 => x"842c728f",
  1636 => x"06535380",
  1637 => x"e2a40880",
  1638 => x"2e9a3872",
  1639 => x"842980e1",
  1640 => x"e4057213",
  1641 => x"81712b70",
  1642 => x"09730806",
  1643 => x"730c5153",
  1644 => x"53b3c704",
  1645 => x"72842980",
  1646 => x"e1e40572",
  1647 => x"1383712b",
  1648 => x"72080772",
  1649 => x"0c535380",
  1650 => x"0b80e2a8",
  1651 => x"0c800b80",
  1652 => x"e2a40c80",
  1653 => x"e49851b4",
  1654 => x"da2d80e3",
  1655 => x"f008ff24",
  1656 => x"feea3880",
  1657 => x"0b80e3f0",
  1658 => x"0c028c05",
  1659 => x"0d0402f8",
  1660 => x"050d80e1",
  1661 => x"e4528f51",
  1662 => x"80727084",
  1663 => x"05540cff",
  1664 => x"11517080",
  1665 => x"25f23802",
  1666 => x"88050d04",
  1667 => x"02f0050d",
  1668 => x"7551b2bf",
  1669 => x"2d70822c",
  1670 => x"fc0680e1",
  1671 => x"e4117210",
  1672 => x"9e067108",
  1673 => x"70722a70",
  1674 => x"83068274",
  1675 => x"2b700974",
  1676 => x"06760c54",
  1677 => x"51565753",
  1678 => x"5153b2b9",
  1679 => x"2d7180e3",
  1680 => x"f00c0290",
  1681 => x"050d0402",
  1682 => x"fc050d72",
  1683 => x"5180710c",
  1684 => x"800b8412",
  1685 => x"0c028405",
  1686 => x"0d0402f0",
  1687 => x"050d7570",
  1688 => x"08841208",
  1689 => x"535353ff",
  1690 => x"5471712e",
  1691 => x"a838b2bf",
  1692 => x"2d841308",
  1693 => x"70842914",
  1694 => x"88117008",
  1695 => x"7081ff06",
  1696 => x"84180881",
  1697 => x"11870684",
  1698 => x"1a0c5351",
  1699 => x"55515151",
  1700 => x"b2b92d71",
  1701 => x"547380e3",
  1702 => x"f00c0290",
  1703 => x"050d0402",
  1704 => x"f8050db2",
  1705 => x"bf2de008",
  1706 => x"708b2a70",
  1707 => x"81065152",
  1708 => x"5270802e",
  1709 => x"a13880e4",
  1710 => x"98087084",
  1711 => x"2980e4a0",
  1712 => x"057381ff",
  1713 => x"06710c51",
  1714 => x"5180e498",
  1715 => x"08811187",
  1716 => x"0680e498",
  1717 => x"0c51800b",
  1718 => x"80e4c00c",
  1719 => x"b2b12db2",
  1720 => x"b92d0288",
  1721 => x"050d0402",
  1722 => x"fc050db2",
  1723 => x"bf2d810b",
  1724 => x"80e4c00c",
  1725 => x"b2b92d80",
  1726 => x"e4c00851",
  1727 => x"70f93802",
  1728 => x"84050d04",
  1729 => x"02fc050d",
  1730 => x"80e49851",
  1731 => x"b4c72db3",
  1732 => x"ee2db59f",
  1733 => x"51b2ad2d",
  1734 => x"0284050d",
  1735 => x"0480e4cc",
  1736 => x"0880e3f0",
  1737 => x"0c0402fc",
  1738 => x"050d810b",
  1739 => x"80e2b00c",
  1740 => x"8151858d",
  1741 => x"2d028405",
  1742 => x"0d0402fc",
  1743 => x"050db6c4",
  1744 => x"04b2c52d",
  1745 => x"80f651b4",
  1746 => x"8c2d80e3",
  1747 => x"f008f238",
  1748 => x"80da51b4",
  1749 => x"8c2d80e3",
  1750 => x"f008e638",
  1751 => x"80e3f008",
  1752 => x"80e2b00c",
  1753 => x"80e3f008",
  1754 => x"51858d2d",
  1755 => x"0284050d",
  1756 => x"0402ec05",
  1757 => x"0d765480",
  1758 => x"52870b88",
  1759 => x"1580f52d",
  1760 => x"56537472",
  1761 => x"248338a0",
  1762 => x"53725183",
  1763 => x"842d8112",
  1764 => x"8b1580f5",
  1765 => x"2d545272",
  1766 => x"7225de38",
  1767 => x"0294050d",
  1768 => x"0402f005",
  1769 => x"0d80e4cc",
  1770 => x"085481f9",
  1771 => x"2d800b80",
  1772 => x"e4d00c73",
  1773 => x"08802e81",
  1774 => x"8938820b",
  1775 => x"80e4840c",
  1776 => x"80e4d008",
  1777 => x"8f0680e4",
  1778 => x"800c7308",
  1779 => x"5271832e",
  1780 => x"96387183",
  1781 => x"26893871",
  1782 => x"812eb038",
  1783 => x"b8ab0471",
  1784 => x"852ea038",
  1785 => x"b8ab0488",
  1786 => x"1480f52d",
  1787 => x"84150880",
  1788 => x"dfa85354",
  1789 => x"5286a02d",
  1790 => x"71842913",
  1791 => x"70085252",
  1792 => x"b8af0473",
  1793 => x"51b6f12d",
  1794 => x"b8ab0480",
  1795 => x"e2ac0888",
  1796 => x"15082c70",
  1797 => x"81065152",
  1798 => x"71802e88",
  1799 => x"3880dfac",
  1800 => x"51b8a804",
  1801 => x"80dfb051",
  1802 => x"86a02d84",
  1803 => x"14085186",
  1804 => x"a02d80e4",
  1805 => x"d0088105",
  1806 => x"80e4d00c",
  1807 => x"8c1454b7",
  1808 => x"b3040290",
  1809 => x"050d0471",
  1810 => x"80e4cc0c",
  1811 => x"b7a12d80",
  1812 => x"e4d008ff",
  1813 => x"0580e4d4",
  1814 => x"0c0402e8",
  1815 => x"050d80e4",
  1816 => x"cc0880e4",
  1817 => x"d8085755",
  1818 => x"80f651b4",
  1819 => x"8c2d80e3",
  1820 => x"f008812a",
  1821 => x"70810651",
  1822 => x"5271802e",
  1823 => x"a438b984",
  1824 => x"04b2c52d",
  1825 => x"80f651b4",
  1826 => x"8c2d80e3",
  1827 => x"f008f238",
  1828 => x"80e2b008",
  1829 => x"81327080",
  1830 => x"e2b00c70",
  1831 => x"5252858d",
  1832 => x"2d800b80",
  1833 => x"e4c40c80",
  1834 => x"0b80e4c8",
  1835 => x"0c80e2b0",
  1836 => x"0883ae38",
  1837 => x"80da51b4",
  1838 => x"8c2d80e3",
  1839 => x"f008802e",
  1840 => x"8c3880e4",
  1841 => x"c4088180",
  1842 => x"0780e4c4",
  1843 => x"0c80d951",
  1844 => x"b48c2d80",
  1845 => x"e3f00880",
  1846 => x"2e8c3880",
  1847 => x"e4c40880",
  1848 => x"c00780e4",
  1849 => x"c40c8194",
  1850 => x"51b48c2d",
  1851 => x"80e3f008",
  1852 => x"802e8b38",
  1853 => x"80e4c408",
  1854 => x"900780e4",
  1855 => x"c40c8191",
  1856 => x"51b48c2d",
  1857 => x"80e3f008",
  1858 => x"802e8b38",
  1859 => x"80e4c408",
  1860 => x"a00780e4",
  1861 => x"c40c81f5",
  1862 => x"51b48c2d",
  1863 => x"80e3f008",
  1864 => x"802e8b38",
  1865 => x"80e4c408",
  1866 => x"810780e4",
  1867 => x"c40c81f2",
  1868 => x"51b48c2d",
  1869 => x"80e3f008",
  1870 => x"802e8b38",
  1871 => x"80e4c408",
  1872 => x"820780e4",
  1873 => x"c40c81eb",
  1874 => x"51b48c2d",
  1875 => x"80e3f008",
  1876 => x"802e8b38",
  1877 => x"80e4c408",
  1878 => x"840780e4",
  1879 => x"c40c81f4",
  1880 => x"51b48c2d",
  1881 => x"80e3f008",
  1882 => x"802e8b38",
  1883 => x"80e4c408",
  1884 => x"880780e4",
  1885 => x"c40c80d8",
  1886 => x"51b48c2d",
  1887 => x"80e3f008",
  1888 => x"802e8c38",
  1889 => x"80e4c808",
  1890 => x"81800780",
  1891 => x"e4c80c92",
  1892 => x"51b48c2d",
  1893 => x"80e3f008",
  1894 => x"802e8c38",
  1895 => x"80e4c808",
  1896 => x"80c00780",
  1897 => x"e4c80c94",
  1898 => x"51b48c2d",
  1899 => x"80e3f008",
  1900 => x"802e8b38",
  1901 => x"80e4c808",
  1902 => x"900780e4",
  1903 => x"c80c9151",
  1904 => x"b48c2d80",
  1905 => x"e3f00880",
  1906 => x"2e8b3880",
  1907 => x"e4c808a0",
  1908 => x"0780e4c8",
  1909 => x"0c9d51b4",
  1910 => x"8c2d80e3",
  1911 => x"f008802e",
  1912 => x"8b3880e4",
  1913 => x"c8088107",
  1914 => x"80e4c80c",
  1915 => x"9b51b48c",
  1916 => x"2d80e3f0",
  1917 => x"08802e8b",
  1918 => x"3880e4c8",
  1919 => x"08820780",
  1920 => x"e4c80c9c",
  1921 => x"51b48c2d",
  1922 => x"80e3f008",
  1923 => x"802e8b38",
  1924 => x"80e4c808",
  1925 => x"840780e4",
  1926 => x"c80ca351",
  1927 => x"b48c2d80",
  1928 => x"e3f00880",
  1929 => x"2e8b3880",
  1930 => x"e4c80888",
  1931 => x"0780e4c8",
  1932 => x"0c9651b4",
  1933 => x"8c2d80e3",
  1934 => x"f008802e",
  1935 => x"843894bf",
  1936 => x"2d9e51b4",
  1937 => x"8c2d80e3",
  1938 => x"f008802e",
  1939 => x"843886ee",
  1940 => x"2d81fd51",
  1941 => x"b48c2d81",
  1942 => x"fa51b48c",
  1943 => x"2d80c2bc",
  1944 => x"0481f551",
  1945 => x"b48c2d80",
  1946 => x"e3f00881",
  1947 => x"2a708106",
  1948 => x"51527180",
  1949 => x"2eb33880",
  1950 => x"e4d40852",
  1951 => x"71802e8a",
  1952 => x"38ff1280",
  1953 => x"e4d40cbd",
  1954 => x"a90480e4",
  1955 => x"d0081080",
  1956 => x"e4d00805",
  1957 => x"70842916",
  1958 => x"51528812",
  1959 => x"08802e89",
  1960 => x"38ff5188",
  1961 => x"12085271",
  1962 => x"2d81f251",
  1963 => x"b48c2d80",
  1964 => x"e3f00881",
  1965 => x"2a708106",
  1966 => x"51527180",
  1967 => x"2eb43880",
  1968 => x"e4d008ff",
  1969 => x"1180e4d4",
  1970 => x"08565353",
  1971 => x"7372258a",
  1972 => x"38811480",
  1973 => x"e4d40cbd",
  1974 => x"f2047210",
  1975 => x"13708429",
  1976 => x"16515288",
  1977 => x"1208802e",
  1978 => x"8938fe51",
  1979 => x"88120852",
  1980 => x"712d81fd",
  1981 => x"51b48c2d",
  1982 => x"80e3f008",
  1983 => x"812a7081",
  1984 => x"06515271",
  1985 => x"802eb138",
  1986 => x"80e4d408",
  1987 => x"802e8a38",
  1988 => x"800b80e4",
  1989 => x"d40cbeb8",
  1990 => x"0480e4d0",
  1991 => x"081080e4",
  1992 => x"d0080570",
  1993 => x"84291651",
  1994 => x"52881208",
  1995 => x"802e8938",
  1996 => x"fd518812",
  1997 => x"0852712d",
  1998 => x"81fa51b4",
  1999 => x"8c2d80e3",
  2000 => x"f008812a",
  2001 => x"70810651",
  2002 => x"5271802e",
  2003 => x"b13880e4",
  2004 => x"d008ff11",
  2005 => x"545280e4",
  2006 => x"d4087325",
  2007 => x"89387280",
  2008 => x"e4d40cbe",
  2009 => x"fe047110",
  2010 => x"12708429",
  2011 => x"16515288",
  2012 => x"1208802e",
  2013 => x"8938fc51",
  2014 => x"88120852",
  2015 => x"712d80e4",
  2016 => x"d4087053",
  2017 => x"5473802e",
  2018 => x"8a388c15",
  2019 => x"ff155555",
  2020 => x"bf850482",
  2021 => x"0b80e484",
  2022 => x"0c718f06",
  2023 => x"80e4800c",
  2024 => x"81eb51b4",
  2025 => x"8c2d80e3",
  2026 => x"f008812a",
  2027 => x"70810651",
  2028 => x"5271802e",
  2029 => x"ad387408",
  2030 => x"852e0981",
  2031 => x"06a43888",
  2032 => x"1580f52d",
  2033 => x"ff055271",
  2034 => x"881681b7",
  2035 => x"2d71982b",
  2036 => x"52718025",
  2037 => x"8838800b",
  2038 => x"881681b7",
  2039 => x"2d7451b6",
  2040 => x"f12d81f4",
  2041 => x"51b48c2d",
  2042 => x"80e3f008",
  2043 => x"812a7081",
  2044 => x"06515271",
  2045 => x"802eb338",
  2046 => x"7408852e",
  2047 => x"098106aa",
  2048 => x"38881580",
  2049 => x"f52d8105",
  2050 => x"52718816",
  2051 => x"81b72d71",
  2052 => x"81ff068b",
  2053 => x"1680f52d",
  2054 => x"54527272",
  2055 => x"27873872",
  2056 => x"881681b7",
  2057 => x"2d7451b6",
  2058 => x"f12d80da",
  2059 => x"51b48c2d",
  2060 => x"80e3f008",
  2061 => x"812a7081",
  2062 => x"06515271",
  2063 => x"802e81b3",
  2064 => x"3880e4cc",
  2065 => x"0880e4d4",
  2066 => x"08555373",
  2067 => x"802e8b38",
  2068 => x"8c13ff15",
  2069 => x"555380c0",
  2070 => x"cb047208",
  2071 => x"5271822e",
  2072 => x"a8387182",
  2073 => x"268a3871",
  2074 => x"812ead38",
  2075 => x"80c1f304",
  2076 => x"71832eb7",
  2077 => x"3871842e",
  2078 => x"09810680",
  2079 => x"f6388813",
  2080 => x"0851b8c7",
  2081 => x"2d80c1f3",
  2082 => x"0480e4d4",
  2083 => x"08518813",
  2084 => x"0852712d",
  2085 => x"80c1f304",
  2086 => x"810b8814",
  2087 => x"082b80e2",
  2088 => x"ac083280",
  2089 => x"e2ac0c80",
  2090 => x"c1c60488",
  2091 => x"1380f52d",
  2092 => x"81058b14",
  2093 => x"80f52d53",
  2094 => x"54717424",
  2095 => x"83388054",
  2096 => x"73881481",
  2097 => x"b72db7a1",
  2098 => x"2d80c1f3",
  2099 => x"04750880",
  2100 => x"2ea43875",
  2101 => x"0851b48c",
  2102 => x"2d80e3f0",
  2103 => x"08810652",
  2104 => x"71802e8c",
  2105 => x"3880e4d4",
  2106 => x"08518416",
  2107 => x"0852712d",
  2108 => x"88165675",
  2109 => x"d8388054",
  2110 => x"800b80e4",
  2111 => x"840c738f",
  2112 => x"0680e480",
  2113 => x"0ca05273",
  2114 => x"80e4d408",
  2115 => x"2e098106",
  2116 => x"993880e4",
  2117 => x"d008ff05",
  2118 => x"74327009",
  2119 => x"81057072",
  2120 => x"079f2a91",
  2121 => x"71315151",
  2122 => x"53537151",
  2123 => x"83842d81",
  2124 => x"14548e74",
  2125 => x"25c23880",
  2126 => x"e2b00852",
  2127 => x"7180e3f0",
  2128 => x"0c029805",
  2129 => x"0d0402f4",
  2130 => x"050dd452",
  2131 => x"81ff720c",
  2132 => x"71085381",
  2133 => x"ff720c72",
  2134 => x"882b83fe",
  2135 => x"80067208",
  2136 => x"7081ff06",
  2137 => x"51525381",
  2138 => x"ff720c72",
  2139 => x"7107882b",
  2140 => x"72087081",
  2141 => x"ff065152",
  2142 => x"5381ff72",
  2143 => x"0c727107",
  2144 => x"882b7208",
  2145 => x"7081ff06",
  2146 => x"720780e3",
  2147 => x"f00c5253",
  2148 => x"028c050d",
  2149 => x"0402f405",
  2150 => x"0d747671",
  2151 => x"81ff06d4",
  2152 => x"0c535380",
  2153 => x"e4dc0885",
  2154 => x"3871892b",
  2155 => x"5271982a",
  2156 => x"d40c7190",
  2157 => x"2a7081ff",
  2158 => x"06d40c51",
  2159 => x"71882a70",
  2160 => x"81ff06d4",
  2161 => x"0c517181",
  2162 => x"ff06d40c",
  2163 => x"72902a70",
  2164 => x"81ff06d4",
  2165 => x"0c51d408",
  2166 => x"7081ff06",
  2167 => x"515182b8",
  2168 => x"bf527081",
  2169 => x"ff2e0981",
  2170 => x"06943881",
  2171 => x"ff0bd40c",
  2172 => x"d4087081",
  2173 => x"ff06ff14",
  2174 => x"54515171",
  2175 => x"e5387080",
  2176 => x"e3f00c02",
  2177 => x"8c050d04",
  2178 => x"02fc050d",
  2179 => x"81c75181",
  2180 => x"ff0bd40c",
  2181 => x"ff115170",
  2182 => x"8025f438",
  2183 => x"0284050d",
  2184 => x"0402f405",
  2185 => x"0d81ff0b",
  2186 => x"d40c9353",
  2187 => x"805287fc",
  2188 => x"80c15180",
  2189 => x"c3952d80",
  2190 => x"e3f0088c",
  2191 => x"3881ff0b",
  2192 => x"d40c8153",
  2193 => x"80c4d204",
  2194 => x"80c4882d",
  2195 => x"ff135372",
  2196 => x"db387280",
  2197 => x"e3f00c02",
  2198 => x"8c050d04",
  2199 => x"02ec050d",
  2200 => x"810b80e4",
  2201 => x"dc0c8454",
  2202 => x"d008708f",
  2203 => x"2a708106",
  2204 => x"51515372",
  2205 => x"f33872d0",
  2206 => x"0c80c488",
  2207 => x"2d80dfb4",
  2208 => x"5186a02d",
  2209 => x"d008708f",
  2210 => x"2a708106",
  2211 => x"51515372",
  2212 => x"f338810b",
  2213 => x"d00cb153",
  2214 => x"805284d4",
  2215 => x"80c05180",
  2216 => x"c3952d80",
  2217 => x"e3f00881",
  2218 => x"2e943872",
  2219 => x"822e80c4",
  2220 => x"38ff1353",
  2221 => x"72e238ff",
  2222 => x"145473ff",
  2223 => x"ab3880c4",
  2224 => x"882d83aa",
  2225 => x"52849c80",
  2226 => x"c85180c3",
  2227 => x"952d80e3",
  2228 => x"f008812e",
  2229 => x"09810694",
  2230 => x"3880c2c6",
  2231 => x"2d80e3f0",
  2232 => x"0883ffff",
  2233 => x"06537283",
  2234 => x"aa2ea338",
  2235 => x"80c4a12d",
  2236 => x"80c68804",
  2237 => x"80dfc051",
  2238 => x"86a02d80",
  2239 => x"5380c7e6",
  2240 => x"0480dfd8",
  2241 => x"5186a02d",
  2242 => x"805480c7",
  2243 => x"b60481ff",
  2244 => x"0bd40cb1",
  2245 => x"5480c488",
  2246 => x"2d8fcf53",
  2247 => x"805287fc",
  2248 => x"80f75180",
  2249 => x"c3952d80",
  2250 => x"e3f00855",
  2251 => x"80e3f008",
  2252 => x"812e0981",
  2253 => x"069e3881",
  2254 => x"ff0bd40c",
  2255 => x"820a5284",
  2256 => x"9c80e951",
  2257 => x"80c3952d",
  2258 => x"80e3f008",
  2259 => x"802e8f38",
  2260 => x"80c4882d",
  2261 => x"ff135372",
  2262 => x"c33880c7",
  2263 => x"a90481ff",
  2264 => x"0bd40c80",
  2265 => x"e3f00852",
  2266 => x"87fc80fa",
  2267 => x"5180c395",
  2268 => x"2d80e3f0",
  2269 => x"08b33881",
  2270 => x"ff0bd40c",
  2271 => x"d4085381",
  2272 => x"ff0bd40c",
  2273 => x"81ff0bd4",
  2274 => x"0c81ff0b",
  2275 => x"d40c81ff",
  2276 => x"0bd40c72",
  2277 => x"862a7081",
  2278 => x"06765651",
  2279 => x"53729738",
  2280 => x"80e3f008",
  2281 => x"5480c7b6",
  2282 => x"0473822e",
  2283 => x"fed338ff",
  2284 => x"145473fe",
  2285 => x"e0387380",
  2286 => x"e4dc0c73",
  2287 => x"8c388152",
  2288 => x"87fc80d0",
  2289 => x"5180c395",
  2290 => x"2d81ff0b",
  2291 => x"d40cd008",
  2292 => x"708f2a70",
  2293 => x"81065151",
  2294 => x"5372f338",
  2295 => x"72d00c81",
  2296 => x"ff0bd40c",
  2297 => x"81537280",
  2298 => x"e3f00c02",
  2299 => x"94050d04",
  2300 => x"02e8050d",
  2301 => x"78558056",
  2302 => x"81ff0bd4",
  2303 => x"0cd00870",
  2304 => x"8f2a7081",
  2305 => x"06515153",
  2306 => x"72f33882",
  2307 => x"810bd00c",
  2308 => x"81ff0bd4",
  2309 => x"0c775287",
  2310 => x"fc80d151",
  2311 => x"80c3952d",
  2312 => x"80dbc6df",
  2313 => x"5480e3f0",
  2314 => x"08802e8c",
  2315 => x"3880dff8",
  2316 => x"5186a02d",
  2317 => x"80c98e04",
  2318 => x"81ff0bd4",
  2319 => x"0cd40870",
  2320 => x"81ff0651",
  2321 => x"537281fe",
  2322 => x"2e098106",
  2323 => x"a03880ff",
  2324 => x"5380c2c6",
  2325 => x"2d80e3f0",
  2326 => x"08757084",
  2327 => x"05570cff",
  2328 => x"13537280",
  2329 => x"25eb3881",
  2330 => x"5680c8f3",
  2331 => x"04ff1454",
  2332 => x"73c63881",
  2333 => x"ff0bd40c",
  2334 => x"81ff0bd4",
  2335 => x"0cd00870",
  2336 => x"8f2a7081",
  2337 => x"06515153",
  2338 => x"72f33872",
  2339 => x"d00c7580",
  2340 => x"e3f00c02",
  2341 => x"98050d04",
  2342 => x"02e8050d",
  2343 => x"77797b58",
  2344 => x"55558053",
  2345 => x"727625a5",
  2346 => x"38747081",
  2347 => x"055680f5",
  2348 => x"2d747081",
  2349 => x"055680f5",
  2350 => x"2d525271",
  2351 => x"712e8738",
  2352 => x"815180c9",
  2353 => x"cf048113",
  2354 => x"5380c9a4",
  2355 => x"04805170",
  2356 => x"80e3f00c",
  2357 => x"0298050d",
  2358 => x"0402ec05",
  2359 => x"0d765574",
  2360 => x"802e80c4",
  2361 => x"389a1580",
  2362 => x"e02d5180",
  2363 => x"d8942d80",
  2364 => x"e3f00880",
  2365 => x"e3f00880",
  2366 => x"eb900c80",
  2367 => x"e3f00854",
  2368 => x"5480eaec",
  2369 => x"08802e9b",
  2370 => x"38941580",
  2371 => x"e02d5180",
  2372 => x"d8942d80",
  2373 => x"e3f00890",
  2374 => x"2b83fff0",
  2375 => x"0a067075",
  2376 => x"07515372",
  2377 => x"80eb900c",
  2378 => x"80eb9008",
  2379 => x"5372802e",
  2380 => x"9e3880ea",
  2381 => x"e408fe14",
  2382 => x"712980ea",
  2383 => x"f8080580",
  2384 => x"eb940c70",
  2385 => x"842b80ea",
  2386 => x"f00c5480",
  2387 => x"cafe0480",
  2388 => x"eafc0880",
  2389 => x"eb900c80",
  2390 => x"eb800880",
  2391 => x"eb940c80",
  2392 => x"eaec0880",
  2393 => x"2e8c3880",
  2394 => x"eae40884",
  2395 => x"2b5380ca",
  2396 => x"f90480eb",
  2397 => x"8408842b",
  2398 => x"537280ea",
  2399 => x"f00c0294",
  2400 => x"050d0402",
  2401 => x"d8050d80",
  2402 => x"0b80eaec",
  2403 => x"0c845480",
  2404 => x"c4dc2d80",
  2405 => x"e3f00880",
  2406 => x"2e993880",
  2407 => x"e4e05280",
  2408 => x"5180c7f0",
  2409 => x"2d80e3f0",
  2410 => x"08802e87",
  2411 => x"38fe5480",
  2412 => x"cbbb04ff",
  2413 => x"14547380",
  2414 => x"24d53873",
  2415 => x"8e3880e0",
  2416 => x"885186a0",
  2417 => x"2d735580",
  2418 => x"d19f0480",
  2419 => x"56810b80",
  2420 => x"eb980c88",
  2421 => x"5380e09c",
  2422 => x"5280e596",
  2423 => x"5180c998",
  2424 => x"2d80e3f0",
  2425 => x"08762e09",
  2426 => x"81068938",
  2427 => x"80e3f008",
  2428 => x"80eb980c",
  2429 => x"885380e0",
  2430 => x"a85280e5",
  2431 => x"b25180c9",
  2432 => x"982d80e3",
  2433 => x"f0088938",
  2434 => x"80e3f008",
  2435 => x"80eb980c",
  2436 => x"80eb9808",
  2437 => x"802e8185",
  2438 => x"3880e8a6",
  2439 => x"0b80f52d",
  2440 => x"80e8a70b",
  2441 => x"80f52d71",
  2442 => x"982b7190",
  2443 => x"2b0780e8",
  2444 => x"a80b80f5",
  2445 => x"2d70882b",
  2446 => x"720780e8",
  2447 => x"a90b80f5",
  2448 => x"2d710780",
  2449 => x"e8de0b80",
  2450 => x"f52d80e8",
  2451 => x"df0b80f5",
  2452 => x"2d71882b",
  2453 => x"07535f54",
  2454 => x"525a5657",
  2455 => x"557381ab",
  2456 => x"aa2e0981",
  2457 => x"06903875",
  2458 => x"5180d7e3",
  2459 => x"2d80e3f0",
  2460 => x"085680cd",
  2461 => x"85047382",
  2462 => x"d4d52e89",
  2463 => x"3880e0b4",
  2464 => x"5180cdd5",
  2465 => x"0480e4e0",
  2466 => x"52755180",
  2467 => x"c7f02d80",
  2468 => x"e3f00855",
  2469 => x"80e3f008",
  2470 => x"802e8483",
  2471 => x"38885380",
  2472 => x"e0a85280",
  2473 => x"e5b25180",
  2474 => x"c9982d80",
  2475 => x"e3f0088b",
  2476 => x"38810b80",
  2477 => x"eaec0c80",
  2478 => x"cddc0488",
  2479 => x"5380e09c",
  2480 => x"5280e596",
  2481 => x"5180c998",
  2482 => x"2d80e3f0",
  2483 => x"08802e8c",
  2484 => x"3880e0c8",
  2485 => x"5186a02d",
  2486 => x"80cebb04",
  2487 => x"80e8de0b",
  2488 => x"80f52d54",
  2489 => x"7380d52e",
  2490 => x"09810680",
  2491 => x"ce3880e8",
  2492 => x"df0b80f5",
  2493 => x"2d547381",
  2494 => x"aa2e0981",
  2495 => x"06bd3880",
  2496 => x"0b80e4e0",
  2497 => x"0b80f52d",
  2498 => x"56547481",
  2499 => x"e92e8338",
  2500 => x"81547481",
  2501 => x"eb2e8c38",
  2502 => x"80557375",
  2503 => x"2e098106",
  2504 => x"82fd3880",
  2505 => x"e4eb0b80",
  2506 => x"f52d5574",
  2507 => x"8e3880e4",
  2508 => x"ec0b80f5",
  2509 => x"2d547382",
  2510 => x"2e873880",
  2511 => x"5580d19f",
  2512 => x"0480e4ed",
  2513 => x"0b80f52d",
  2514 => x"7080eae4",
  2515 => x"0cff0580",
  2516 => x"eae80c80",
  2517 => x"e4ee0b80",
  2518 => x"f52d80e4",
  2519 => x"ef0b80f5",
  2520 => x"2d587605",
  2521 => x"77828029",
  2522 => x"057080ea",
  2523 => x"f40c80e4",
  2524 => x"f00b80f5",
  2525 => x"2d7080eb",
  2526 => x"880c80ea",
  2527 => x"ec085957",
  2528 => x"5876802e",
  2529 => x"81b93888",
  2530 => x"5380e0a8",
  2531 => x"5280e5b2",
  2532 => x"5180c998",
  2533 => x"2d80e3f0",
  2534 => x"08828438",
  2535 => x"80eae408",
  2536 => x"70842b80",
  2537 => x"eaf00c70",
  2538 => x"80eb840c",
  2539 => x"80e5850b",
  2540 => x"80f52d80",
  2541 => x"e5840b80",
  2542 => x"f52d7182",
  2543 => x"80290580",
  2544 => x"e5860b80",
  2545 => x"f52d7084",
  2546 => x"80802912",
  2547 => x"80e5870b",
  2548 => x"80f52d70",
  2549 => x"81800a29",
  2550 => x"127080eb",
  2551 => x"8c0c80eb",
  2552 => x"88087129",
  2553 => x"80eaf408",
  2554 => x"057080ea",
  2555 => x"f80c80e5",
  2556 => x"8d0b80f5",
  2557 => x"2d80e58c",
  2558 => x"0b80f52d",
  2559 => x"71828029",
  2560 => x"0580e58e",
  2561 => x"0b80f52d",
  2562 => x"70848080",
  2563 => x"291280e5",
  2564 => x"8f0b80f5",
  2565 => x"2d70982b",
  2566 => x"81f00a06",
  2567 => x"72057080",
  2568 => x"eafc0cfe",
  2569 => x"117e2977",
  2570 => x"0580eb80",
  2571 => x"0c525952",
  2572 => x"43545e51",
  2573 => x"5259525d",
  2574 => x"57595780",
  2575 => x"d1970480",
  2576 => x"e4f20b80",
  2577 => x"f52d80e4",
  2578 => x"f10b80f5",
  2579 => x"2d718280",
  2580 => x"29057080",
  2581 => x"eaf00c70",
  2582 => x"a02983ff",
  2583 => x"0570892a",
  2584 => x"7080eb84",
  2585 => x"0c80e4f7",
  2586 => x"0b80f52d",
  2587 => x"80e4f60b",
  2588 => x"80f52d71",
  2589 => x"82802905",
  2590 => x"7080eb8c",
  2591 => x"0c7b7129",
  2592 => x"1e7080eb",
  2593 => x"800c7d80",
  2594 => x"eafc0c73",
  2595 => x"0580eaf8",
  2596 => x"0c555e51",
  2597 => x"51555580",
  2598 => x"5180c9d9",
  2599 => x"2d815574",
  2600 => x"80e3f00c",
  2601 => x"02a8050d",
  2602 => x"0402ec05",
  2603 => x"0d767087",
  2604 => x"2c7180ff",
  2605 => x"06555654",
  2606 => x"80eaec08",
  2607 => x"8a387388",
  2608 => x"2c7481ff",
  2609 => x"06545580",
  2610 => x"e4e05280",
  2611 => x"eaf40815",
  2612 => x"5180c7f0",
  2613 => x"2d80e3f0",
  2614 => x"085480e3",
  2615 => x"f008802e",
  2616 => x"bb3880ea",
  2617 => x"ec08802e",
  2618 => x"9c387284",
  2619 => x"2980e4e0",
  2620 => x"05700852",
  2621 => x"5380d7e3",
  2622 => x"2d80e3f0",
  2623 => x"08f00a06",
  2624 => x"5380d29a",
  2625 => x"04721080",
  2626 => x"e4e00570",
  2627 => x"80e02d52",
  2628 => x"5380d894",
  2629 => x"2d80e3f0",
  2630 => x"08537254",
  2631 => x"7380e3f0",
  2632 => x"0c029405",
  2633 => x"0d0402e0",
  2634 => x"050d7970",
  2635 => x"842c80eb",
  2636 => x"94080571",
  2637 => x"8f065255",
  2638 => x"53728b38",
  2639 => x"80e4e052",
  2640 => x"735180c7",
  2641 => x"f02d72a0",
  2642 => x"2980e4e0",
  2643 => x"05548074",
  2644 => x"80f52d56",
  2645 => x"5374732e",
  2646 => x"83388153",
  2647 => x"7481e52e",
  2648 => x"81f53881",
  2649 => x"70740654",
  2650 => x"5872802e",
  2651 => x"81e9388b",
  2652 => x"1480f52d",
  2653 => x"70832a79",
  2654 => x"06585676",
  2655 => x"9c3880e2",
  2656 => x"b4085372",
  2657 => x"89387280",
  2658 => x"e8e00b81",
  2659 => x"b72d7680",
  2660 => x"e2b40c73",
  2661 => x"5380d4d9",
  2662 => x"04758f2e",
  2663 => x"09810681",
  2664 => x"b638749f",
  2665 => x"068d2980",
  2666 => x"e8d31151",
  2667 => x"53811480",
  2668 => x"f52d7370",
  2669 => x"81055581",
  2670 => x"b72d8314",
  2671 => x"80f52d73",
  2672 => x"70810555",
  2673 => x"81b72d85",
  2674 => x"1480f52d",
  2675 => x"73708105",
  2676 => x"5581b72d",
  2677 => x"871480f5",
  2678 => x"2d737081",
  2679 => x"055581b7",
  2680 => x"2d891480",
  2681 => x"f52d7370",
  2682 => x"81055581",
  2683 => x"b72d8e14",
  2684 => x"80f52d73",
  2685 => x"70810555",
  2686 => x"81b72d90",
  2687 => x"1480f52d",
  2688 => x"73708105",
  2689 => x"5581b72d",
  2690 => x"921480f5",
  2691 => x"2d737081",
  2692 => x"055581b7",
  2693 => x"2d941480",
  2694 => x"f52d7370",
  2695 => x"81055581",
  2696 => x"b72d9614",
  2697 => x"80f52d73",
  2698 => x"70810555",
  2699 => x"81b72d98",
  2700 => x"1480f52d",
  2701 => x"73708105",
  2702 => x"5581b72d",
  2703 => x"9c1480f5",
  2704 => x"2d737081",
  2705 => x"055581b7",
  2706 => x"2d9e1480",
  2707 => x"f52d7381",
  2708 => x"b72d7780",
  2709 => x"e2b40c80",
  2710 => x"537280e3",
  2711 => x"f00c02a0",
  2712 => x"050d0402",
  2713 => x"cc050d7e",
  2714 => x"605e5a80",
  2715 => x"0b80eb90",
  2716 => x"0880eb94",
  2717 => x"08595c56",
  2718 => x"805880ea",
  2719 => x"f008782e",
  2720 => x"81be3877",
  2721 => x"8f06a017",
  2722 => x"57547392",
  2723 => x"3880e4e0",
  2724 => x"52765181",
  2725 => x"175780c7",
  2726 => x"f02d80e4",
  2727 => x"e0568076",
  2728 => x"80f52d56",
  2729 => x"5474742e",
  2730 => x"83388154",
  2731 => x"7481e52e",
  2732 => x"81823881",
  2733 => x"70750655",
  2734 => x"5c73802e",
  2735 => x"80f6388b",
  2736 => x"1680f52d",
  2737 => x"98065978",
  2738 => x"80ea388b",
  2739 => x"537c5275",
  2740 => x"5180c998",
  2741 => x"2d80e3f0",
  2742 => x"0880d938",
  2743 => x"9c160851",
  2744 => x"80d7e32d",
  2745 => x"80e3f008",
  2746 => x"841b0c9a",
  2747 => x"1680e02d",
  2748 => x"5180d894",
  2749 => x"2d80e3f0",
  2750 => x"0880e3f0",
  2751 => x"08881c0c",
  2752 => x"80e3f008",
  2753 => x"555580ea",
  2754 => x"ec08802e",
  2755 => x"9a389416",
  2756 => x"80e02d51",
  2757 => x"80d8942d",
  2758 => x"80e3f008",
  2759 => x"902b83ff",
  2760 => x"f00a0670",
  2761 => x"16515473",
  2762 => x"881b0c78",
  2763 => x"7a0c7b54",
  2764 => x"80d6fe04",
  2765 => x"81185880",
  2766 => x"eaf00878",
  2767 => x"26fec438",
  2768 => x"80eaec08",
  2769 => x"802eb538",
  2770 => x"7a5180d1",
  2771 => x"a92d80e3",
  2772 => x"f00880e3",
  2773 => x"f00880ff",
  2774 => x"fffff806",
  2775 => x"555b7380",
  2776 => x"fffffff8",
  2777 => x"2e963880",
  2778 => x"e3f008fe",
  2779 => x"0580eae4",
  2780 => x"082980ea",
  2781 => x"f8080557",
  2782 => x"80d4f804",
  2783 => x"80547380",
  2784 => x"e3f00c02",
  2785 => x"b4050d04",
  2786 => x"02f4050d",
  2787 => x"74700881",
  2788 => x"05710c70",
  2789 => x"0880eae8",
  2790 => x"08065353",
  2791 => x"71903888",
  2792 => x"13085180",
  2793 => x"d1a92d80",
  2794 => x"e3f00888",
  2795 => x"140c810b",
  2796 => x"80e3f00c",
  2797 => x"028c050d",
  2798 => x"0402f005",
  2799 => x"0d758811",
  2800 => x"08fe0580",
  2801 => x"eae40829",
  2802 => x"80eaf808",
  2803 => x"11720880",
  2804 => x"eae80806",
  2805 => x"05795553",
  2806 => x"545480c7",
  2807 => x"f02d0290",
  2808 => x"050d0402",
  2809 => x"f4050d74",
  2810 => x"70882a83",
  2811 => x"fe800670",
  2812 => x"72982a07",
  2813 => x"72882b87",
  2814 => x"fc808006",
  2815 => x"73982b81",
  2816 => x"f00a0671",
  2817 => x"73070780",
  2818 => x"e3f00c56",
  2819 => x"51535102",
  2820 => x"8c050d04",
  2821 => x"02f8050d",
  2822 => x"028e0580",
  2823 => x"f52d7488",
  2824 => x"2b077083",
  2825 => x"ffff0680",
  2826 => x"e3f00c51",
  2827 => x"0288050d",
  2828 => x"0402f405",
  2829 => x"0d747678",
  2830 => x"53545280",
  2831 => x"71259738",
  2832 => x"72708105",
  2833 => x"5480f52d",
  2834 => x"72708105",
  2835 => x"5481b72d",
  2836 => x"ff115170",
  2837 => x"eb388072",
  2838 => x"81b72d02",
  2839 => x"8c050d04",
  2840 => x"02e8050d",
  2841 => x"77568070",
  2842 => x"56547376",
  2843 => x"24b73880",
  2844 => x"eaf00874",
  2845 => x"2eaf3873",
  2846 => x"5180d2a6",
  2847 => x"2d80e3f0",
  2848 => x"0880e3f0",
  2849 => x"08098105",
  2850 => x"7080e3f0",
  2851 => x"08079f2a",
  2852 => x"77058117",
  2853 => x"57575353",
  2854 => x"74762489",
  2855 => x"3880eaf0",
  2856 => x"087426d3",
  2857 => x"387280e3",
  2858 => x"f00c0298",
  2859 => x"050d0402",
  2860 => x"f0050d80",
  2861 => x"e3ec0816",
  2862 => x"5180d8e0",
  2863 => x"2d80e3f0",
  2864 => x"08802ea0",
  2865 => x"388b5380",
  2866 => x"e3f00852",
  2867 => x"80e8e051",
  2868 => x"80d8b12d",
  2869 => x"80eb9c08",
  2870 => x"5473802e",
  2871 => x"873880e8",
  2872 => x"e051732d",
  2873 => x"0290050d",
  2874 => x"0402dc05",
  2875 => x"0d80705a",
  2876 => x"557480e3",
  2877 => x"ec0825b5",
  2878 => x"3880eaf0",
  2879 => x"08752ead",
  2880 => x"38785180",
  2881 => x"d2a62d80",
  2882 => x"e3f00809",
  2883 => x"81057080",
  2884 => x"e3f00807",
  2885 => x"9f2a7605",
  2886 => x"811b5b56",
  2887 => x"547480e3",
  2888 => x"ec082589",
  2889 => x"3880eaf0",
  2890 => x"087926d5",
  2891 => x"38805578",
  2892 => x"80eaf008",
  2893 => x"2781e438",
  2894 => x"785180d2",
  2895 => x"a62d80e3",
  2896 => x"f008802e",
  2897 => x"81b43880",
  2898 => x"e3f0088b",
  2899 => x"0580f52d",
  2900 => x"70842a70",
  2901 => x"81067710",
  2902 => x"78842b80",
  2903 => x"e8e00b80",
  2904 => x"f52d5c5c",
  2905 => x"53515556",
  2906 => x"73802e80",
  2907 => x"ce387416",
  2908 => x"822b80dc",
  2909 => x"bf0b80e2",
  2910 => x"c0120c54",
  2911 => x"77753110",
  2912 => x"80eba011",
  2913 => x"55569074",
  2914 => x"70810556",
  2915 => x"81b72da0",
  2916 => x"7481b72d",
  2917 => x"7681ff06",
  2918 => x"81165854",
  2919 => x"73802e8b",
  2920 => x"389c5380",
  2921 => x"e8e05280",
  2922 => x"dbb2048b",
  2923 => x"5380e3f0",
  2924 => x"085280eb",
  2925 => x"a2165180",
  2926 => x"dbf00474",
  2927 => x"16822b80",
  2928 => x"d9af0b80",
  2929 => x"e2c0120c",
  2930 => x"547681ff",
  2931 => x"06811658",
  2932 => x"5473802e",
  2933 => x"8b389c53",
  2934 => x"80e8e052",
  2935 => x"80dbe704",
  2936 => x"8b5380e3",
  2937 => x"f0085277",
  2938 => x"75311080",
  2939 => x"eba00551",
  2940 => x"765580d8",
  2941 => x"b12d80dc",
  2942 => x"8f047490",
  2943 => x"29753170",
  2944 => x"1080eba0",
  2945 => x"05515480",
  2946 => x"e3f00874",
  2947 => x"81b72d81",
  2948 => x"1959748b",
  2949 => x"24a43880",
  2950 => x"daaf0474",
  2951 => x"90297531",
  2952 => x"701080eb",
  2953 => x"a0058c77",
  2954 => x"31575154",
  2955 => x"807481b7",
  2956 => x"2d9e14ff",
  2957 => x"16565474",
  2958 => x"f33802a4",
  2959 => x"050d0402",
  2960 => x"fc050d80",
  2961 => x"e3ec0813",
  2962 => x"5180d8e0",
  2963 => x"2d80e3f0",
  2964 => x"08802e8a",
  2965 => x"3880e3f0",
  2966 => x"085180c9",
  2967 => x"d92d800b",
  2968 => x"80e3ec0c",
  2969 => x"80d9e92d",
  2970 => x"b7a12d02",
  2971 => x"84050d04",
  2972 => x"02fc050d",
  2973 => x"725170fd",
  2974 => x"2eb23870",
  2975 => x"fd248b38",
  2976 => x"70fc2e80",
  2977 => x"d03880dd",
  2978 => x"df0470fe",
  2979 => x"2eb93870",
  2980 => x"ff2e0981",
  2981 => x"0680c838",
  2982 => x"80e3ec08",
  2983 => x"5170802e",
  2984 => x"be38ff11",
  2985 => x"80e3ec0c",
  2986 => x"80dddf04",
  2987 => x"80e3ec08",
  2988 => x"f0057080",
  2989 => x"e3ec0c51",
  2990 => x"708025a3",
  2991 => x"38800b80",
  2992 => x"e3ec0c80",
  2993 => x"dddf0480",
  2994 => x"e3ec0881",
  2995 => x"0580e3ec",
  2996 => x"0c80dddf",
  2997 => x"0480e3ec",
  2998 => x"08900580",
  2999 => x"e3ec0c80",
  3000 => x"d9e92db7",
  3001 => x"a12d0284",
  3002 => x"050d0402",
  3003 => x"fc050d80",
  3004 => x"0b80e3ec",
  3005 => x"0c80d9e9",
  3006 => x"2db69d2d",
  3007 => x"80e3f008",
  3008 => x"80e3dc0c",
  3009 => x"80e2b851",
  3010 => x"b8c72d02",
  3011 => x"84050d04",
  3012 => x"7180eb9c",
  3013 => x"0c040000",
  3014 => x"00ffffff",
  3015 => x"ff00ffff",
  3016 => x"ffff00ff",
  3017 => x"ffffff00",
  3018 => x"52657365",
  3019 => x"74204e45",
  3020 => x"53000000",
  3021 => x"5363616e",
  3022 => x"6c696e65",
  3023 => x"73000000",
  3024 => x"48513258",
  3025 => x"2046696c",
  3026 => x"74657200",
  3027 => x"50312053",
  3028 => x"656c6563",
  3029 => x"74000000",
  3030 => x"50312053",
  3031 => x"74617274",
  3032 => x"00000000",
  3033 => x"4c6f6164",
  3034 => x"20524f4d",
  3035 => x"20100000",
  3036 => x"45786974",
  3037 => x"00000000",
  3038 => x"524f4d20",
  3039 => x"6c6f6164",
  3040 => x"696e6720",
  3041 => x"6661696c",
  3042 => x"65640000",
  3043 => x"4f4b0000",
  3044 => x"496e6974",
  3045 => x"69616c69",
  3046 => x"7a696e67",
  3047 => x"20534420",
  3048 => x"63617264",
  3049 => x"0a000000",
  3050 => x"16200000",
  3051 => x"14200000",
  3052 => x"15200000",
  3053 => x"53442069",
  3054 => x"6e69742e",
  3055 => x"2e2e0a00",
  3056 => x"53442063",
  3057 => x"61726420",
  3058 => x"72657365",
  3059 => x"74206661",
  3060 => x"696c6564",
  3061 => x"210a0000",
  3062 => x"53444843",
  3063 => x"20657272",
  3064 => x"6f72210a",
  3065 => x"00000000",
  3066 => x"57726974",
  3067 => x"65206661",
  3068 => x"696c6564",
  3069 => x"0a000000",
  3070 => x"52656164",
  3071 => x"20666169",
  3072 => x"6c65640a",
  3073 => x"00000000",
  3074 => x"43617264",
  3075 => x"20696e69",
  3076 => x"74206661",
  3077 => x"696c6564",
  3078 => x"0a000000",
  3079 => x"46415431",
  3080 => x"36202020",
  3081 => x"00000000",
  3082 => x"46415433",
  3083 => x"32202020",
  3084 => x"00000000",
  3085 => x"4e6f2070",
  3086 => x"61727469",
  3087 => x"74696f6e",
  3088 => x"20736967",
  3089 => x"0a000000",
  3090 => x"42616420",
  3091 => x"70617274",
  3092 => x"0a000000",
  3093 => x"4261636b",
  3094 => x"00000000",
  3095 => x"00000002",
  3096 => x"00000002",
  3097 => x"00002f28",
  3098 => x"0000035a",
  3099 => x"00000001",
  3100 => x"00002f34",
  3101 => x"00000000",
  3102 => x"00000001",
  3103 => x"00002f40",
  3104 => x"00000001",
  3105 => x"00000002",
  3106 => x"00002f4c",
  3107 => x"0000036e",
  3108 => x"00000002",
  3109 => x"00002f58",
  3110 => x"00000a3f",
  3111 => x"00000002",
  3112 => x"00002f64",
  3113 => x"00002eeb",
  3114 => x"00000002",
  3115 => x"00002f70",
  3116 => x"00001b3a",
  3117 => x"00000000",
  3118 => x"00000000",
  3119 => x"00000000",
  3120 => x"00000004",
  3121 => x"00002f78",
  3122 => x"000030c0",
  3123 => x"00000004",
  3124 => x"00002f8c",
  3125 => x"00003060",
  3126 => x"00000000",
  3127 => x"00000000",
  3128 => x"00000000",
  3129 => x"00000000",
  3130 => x"00000000",
  3131 => x"00000000",
  3132 => x"00000000",
  3133 => x"00000000",
  3134 => x"00000000",
  3135 => x"00000000",
  3136 => x"00000000",
  3137 => x"00000000",
  3138 => x"00000000",
  3139 => x"00000000",
  3140 => x"00000000",
  3141 => x"00000000",
  3142 => x"00000000",
  3143 => x"00000000",
  3144 => x"00000000",
  3145 => x"00000000",
  3146 => x"00000000",
  3147 => x"00000000",
  3148 => x"00000000",
  3149 => x"00000000",
  3150 => x"00000002",
  3151 => x"000035a0",
  3152 => x"00002caf",
  3153 => x"00000002",
  3154 => x"000035be",
  3155 => x"00002caf",
  3156 => x"00000002",
  3157 => x"000035dc",
  3158 => x"00002caf",
  3159 => x"00000002",
  3160 => x"000035fa",
  3161 => x"00002caf",
  3162 => x"00000002",
  3163 => x"00003618",
  3164 => x"00002caf",
  3165 => x"00000002",
  3166 => x"00003636",
  3167 => x"00002caf",
  3168 => x"00000002",
  3169 => x"00003654",
  3170 => x"00002caf",
  3171 => x"00000002",
  3172 => x"00003672",
  3173 => x"00002caf",
  3174 => x"00000002",
  3175 => x"00003690",
  3176 => x"00002caf",
  3177 => x"00000002",
  3178 => x"000036ae",
  3179 => x"00002caf",
  3180 => x"00000002",
  3181 => x"000036cc",
  3182 => x"00002caf",
  3183 => x"00000002",
  3184 => x"000036ea",
  3185 => x"00002caf",
  3186 => x"00000002",
  3187 => x"00003708",
  3188 => x"00002caf",
  3189 => x"00000004",
  3190 => x"00003054",
  3191 => x"00000000",
  3192 => x"00000000",
  3193 => x"00000000",
  3194 => x"00002e70",
  3195 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

