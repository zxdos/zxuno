-------------------------------------------------------------------------------
--
-- $Id: T80_Reg-c.vhd,v 1.1 2006/01/03 08:23:24 arnim Exp $
--
-------------------------------------------------------------------------------

configuration T80_Reg_rtl_c0 of T80_Reg is

  for rtl
  end for;

end T80_Reg_rtl_c0;
